library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use WORK.constants.all;

entity LUT_ROM is
	generic (
		N : integer := N_WRF;
		F : integer := F_WRF;
		M : integer := M_WRF
	);
	port(
		Clk : in std_logic;
		addr1, addr2 : in std_logic_vector(integer(ceil(log2(real(3*N + M) + real(1))))-1 downto 0); -- address 
		en   : in std_logic_vector(F-1 downto 0); -- ROM Enable, for additiona
		dout1, dout2 : out std_logic_vector(integer(ceil(log2(real(2*N*F + M) + real(1))))-1 downto 0)
	);
end entity;

architecture beh of LUT_ROM is 
begin


    -- Output port #1
    process(Clk, addr1, en)
        variable en_addr : std_logic_vector(8+5-1 downto 0);
    begin
        en_addr := en & addr1;
        if (rising_edge(Clk)) then 
            case (en_addr) is
        -- block #1

        -- 3*N registers for IN/LOC/OUT registers
                when "1000000000000" =>
                    dout1 <= "00000000";
                when "1000000000001" =>
                    dout1 <= "00000001";
                when "1000000000010" =>
                    dout1 <= "00000010";
                when "1000000000011" =>
                    dout1 <= "00000011";
                when "1000000000100" =>
                    dout1 <= "00000100";
                when "1000000000101" =>
                    dout1 <= "00000101";
                when "1000000000110" =>
                    dout1 <= "00000110";
                when "1000000000111" =>
                    dout1 <= "00000111";
                when "1000000001000" =>
                    dout1 <= "00001000";
                when "1000000001001" =>
                    dout1 <= "00001001";
                when "1000000001010" =>
                    dout1 <= "00001010";
                when "1000000001011" =>
                    dout1 <= "00001011";
                when "1000000001100" =>
                    dout1 <= "00001100";
                when "1000000001101" =>
                    dout1 <= "00001101";
                when "1000000001110" =>
                    dout1 <= "00001110";
                when "1000000001111" =>
                    dout1 <= "00001111";
                when "1000000010000" =>
                    dout1 <= "00010000";
                when "1000000010001" =>
                    dout1 <= "00010001";
                when "1000000010010" =>
                    dout1 <= "00010010";
                when "1000000010011" =>
                    dout1 <= "00010011";
                when "1000000010100" =>
                    dout1 <= "00010100";
                when "1000000010101" =>
                    dout1 <= "00010101";
                when "1000000010110" =>
                    dout1 <= "00010110";
                when "1000000010111" =>
                    dout1 <= "00010111";

    -- M global registers
                when "1000000011000" =>
                    dout1 <= "10000000";
                when "1000000011001" =>
                    dout1 <= "10000001";
                when "1000000011010" =>
                    dout1 <= "10000010";

        -- block #2

        -- 3*N registers for IN/LOC/OUT registers
                when "0100000000000" =>
                    dout1 <= "00010000";
                when "0100000000001" =>
                    dout1 <= "00010001";
                when "0100000000010" =>
                    dout1 <= "00010010";
                when "0100000000011" =>
                    dout1 <= "00010011";
                when "0100000000100" =>
                    dout1 <= "00010100";
                when "0100000000101" =>
                    dout1 <= "00010101";
                when "0100000000110" =>
                    dout1 <= "00010110";
                when "0100000000111" =>
                    dout1 <= "00010111";
                when "0100000001000" =>
                    dout1 <= "00011000";
                when "0100000001001" =>
                    dout1 <= "00011001";
                when "0100000001010" =>
                    dout1 <= "00011010";
                when "0100000001011" =>
                    dout1 <= "00011011";
                when "0100000001100" =>
                    dout1 <= "00011100";
                when "0100000001101" =>
                    dout1 <= "00011101";
                when "0100000001110" =>
                    dout1 <= "00011110";
                when "0100000001111" =>
                    dout1 <= "00011111";
                when "0100000010000" =>
                    dout1 <= "00100000";
                when "0100000010001" =>
                    dout1 <= "00100001";
                when "0100000010010" =>
                    dout1 <= "00100010";
                when "0100000010011" =>
                    dout1 <= "00100011";
                when "0100000010100" =>
                    dout1 <= "00100100";
                when "0100000010101" =>
                    dout1 <= "00100101";
                when "0100000010110" =>
                    dout1 <= "00100110";
                when "0100000010111" =>
                    dout1 <= "00100111";

    -- M global registers
                when "0100000011000" =>
                    dout1 <= "10000000";
                when "0100000011001" =>
                    dout1 <= "10000001";
                when "0100000011010" =>
                    dout1 <= "10000010";

        -- block #3

        -- 3*N registers for IN/LOC/OUT registers
                when "0010000000000" =>
                    dout1 <= "00100000";
                when "0010000000001" =>
                    dout1 <= "00100001";
                when "0010000000010" =>
                    dout1 <= "00100010";
                when "0010000000011" =>
                    dout1 <= "00100011";
                when "0010000000100" =>
                    dout1 <= "00100100";
                when "0010000000101" =>
                    dout1 <= "00100101";
                when "0010000000110" =>
                    dout1 <= "00100110";
                when "0010000000111" =>
                    dout1 <= "00100111";
                when "0010000001000" =>
                    dout1 <= "00101000";
                when "0010000001001" =>
                    dout1 <= "00101001";
                when "0010000001010" =>
                    dout1 <= "00101010";
                when "0010000001011" =>
                    dout1 <= "00101011";
                when "0010000001100" =>
                    dout1 <= "00101100";
                when "0010000001101" =>
                    dout1 <= "00101101";
                when "0010000001110" =>
                    dout1 <= "00101110";
                when "0010000001111" =>
                    dout1 <= "00101111";
                when "0010000010000" =>
                    dout1 <= "00110000";
                when "0010000010001" =>
                    dout1 <= "00110001";
                when "0010000010010" =>
                    dout1 <= "00110010";
                when "0010000010011" =>
                    dout1 <= "00110011";
                when "0010000010100" =>
                    dout1 <= "00110100";
                when "0010000010101" =>
                    dout1 <= "00110101";
                when "0010000010110" =>
                    dout1 <= "00110110";
                when "0010000010111" =>
                    dout1 <= "00110111";

    -- M global registers
                when "0010000011000" =>
                    dout1 <= "10000000";
                when "0010000011001" =>
                    dout1 <= "10000001";
                when "0010000011010" =>
                    dout1 <= "10000010";

        -- block #4

        -- 3*N registers for IN/LOC/OUT registers
                when "0001000000000" =>
                    dout1 <= "00110000";
                when "0001000000001" =>
                    dout1 <= "00110001";
                when "0001000000010" =>
                    dout1 <= "00110010";
                when "0001000000011" =>
                    dout1 <= "00110011";
                when "0001000000100" =>
                    dout1 <= "00110100";
                when "0001000000101" =>
                    dout1 <= "00110101";
                when "0001000000110" =>
                    dout1 <= "00110110";
                when "0001000000111" =>
                    dout1 <= "00110111";
                when "0001000001000" =>
                    dout1 <= "00111000";
                when "0001000001001" =>
                    dout1 <= "00111001";
                when "0001000001010" =>
                    dout1 <= "00111010";
                when "0001000001011" =>
                    dout1 <= "00111011";
                when "0001000001100" =>
                    dout1 <= "00111100";
                when "0001000001101" =>
                    dout1 <= "00111101";
                when "0001000001110" =>
                    dout1 <= "00111110";
                when "0001000001111" =>
                    dout1 <= "00111111";
                when "0001000010000" =>
                    dout1 <= "01000000";
                when "0001000010001" =>
                    dout1 <= "01000001";
                when "0001000010010" =>
                    dout1 <= "01000010";
                when "0001000010011" =>
                    dout1 <= "01000011";
                when "0001000010100" =>
                    dout1 <= "01000100";
                when "0001000010101" =>
                    dout1 <= "01000101";
                when "0001000010110" =>
                    dout1 <= "01000110";
                when "0001000010111" =>
                    dout1 <= "01000111";

    -- M global registers
                when "0001000011000" =>
                    dout1 <= "10000000";
                when "0001000011001" =>
                    dout1 <= "10000001";
                when "0001000011010" =>
                    dout1 <= "10000010";

        -- block #5

        -- 3*N registers for IN/LOC/OUT registers
                when "0000100000000" =>
                    dout1 <= "01000000";
                when "0000100000001" =>
                    dout1 <= "01000001";
                when "0000100000010" =>
                    dout1 <= "01000010";
                when "0000100000011" =>
                    dout1 <= "01000011";
                when "0000100000100" =>
                    dout1 <= "01000100";
                when "0000100000101" =>
                    dout1 <= "01000101";
                when "0000100000110" =>
                    dout1 <= "01000110";
                when "0000100000111" =>
                    dout1 <= "01000111";
                when "0000100001000" =>
                    dout1 <= "01001000";
                when "0000100001001" =>
                    dout1 <= "01001001";
                when "0000100001010" =>
                    dout1 <= "01001010";
                when "0000100001011" =>
                    dout1 <= "01001011";
                when "0000100001100" =>
                    dout1 <= "01001100";
                when "0000100001101" =>
                    dout1 <= "01001101";
                when "0000100001110" =>
                    dout1 <= "01001110";
                when "0000100001111" =>
                    dout1 <= "01001111";
                when "0000100010000" =>
                    dout1 <= "01010000";
                when "0000100010001" =>
                    dout1 <= "01010001";
                when "0000100010010" =>
                    dout1 <= "01010010";
                when "0000100010011" =>
                    dout1 <= "01010011";
                when "0000100010100" =>
                    dout1 <= "01010100";
                when "0000100010101" =>
                    dout1 <= "01010101";
                when "0000100010110" =>
                    dout1 <= "01010110";
                when "0000100010111" =>
                    dout1 <= "01010111";

    -- M global registers
                when "0000100011000" =>
                    dout1 <= "10000000";
                when "0000100011001" =>
                    dout1 <= "10000001";
                when "0000100011010" =>
                    dout1 <= "10000010";

        -- block #6

        -- 3*N registers for IN/LOC/OUT registers
                when "0000010000000" =>
                    dout1 <= "01010000";
                when "0000010000001" =>
                    dout1 <= "01010001";
                when "0000010000010" =>
                    dout1 <= "01010010";
                when "0000010000011" =>
                    dout1 <= "01010011";
                when "0000010000100" =>
                    dout1 <= "01010100";
                when "0000010000101" =>
                    dout1 <= "01010101";
                when "0000010000110" =>
                    dout1 <= "01010110";
                when "0000010000111" =>
                    dout1 <= "01010111";
                when "0000010001000" =>
                    dout1 <= "01011000";
                when "0000010001001" =>
                    dout1 <= "01011001";
                when "0000010001010" =>
                    dout1 <= "01011010";
                when "0000010001011" =>
                    dout1 <= "01011011";
                when "0000010001100" =>
                    dout1 <= "01011100";
                when "0000010001101" =>
                    dout1 <= "01011101";
                when "0000010001110" =>
                    dout1 <= "01011110";
                when "0000010001111" =>
                    dout1 <= "01011111";
                when "0000010010000" =>
                    dout1 <= "01100000";
                when "0000010010001" =>
                    dout1 <= "01100001";
                when "0000010010010" =>
                    dout1 <= "01100010";
                when "0000010010011" =>
                    dout1 <= "01100011";
                when "0000010010100" =>
                    dout1 <= "01100100";
                when "0000010010101" =>
                    dout1 <= "01100101";
                when "0000010010110" =>
                    dout1 <= "01100110";
                when "0000010010111" =>
                    dout1 <= "01100111";

    -- M global registers
                when "0000010011000" =>
                    dout1 <= "10000000";
                when "0000010011001" =>
                    dout1 <= "10000001";
                when "0000010011010" =>
                    dout1 <= "10000010";

        -- block #7

        -- 3*N registers for IN/LOC/OUT registers
                when "0000001000000" =>
                    dout1 <= "01100000";
                when "0000001000001" =>
                    dout1 <= "01100001";
                when "0000001000010" =>
                    dout1 <= "01100010";
                when "0000001000011" =>
                    dout1 <= "01100011";
                when "0000001000100" =>
                    dout1 <= "01100100";
                when "0000001000101" =>
                    dout1 <= "01100101";
                when "0000001000110" =>
                    dout1 <= "01100110";
                when "0000001000111" =>
                    dout1 <= "01100111";
                when "0000001001000" =>
                    dout1 <= "01101000";
                when "0000001001001" =>
                    dout1 <= "01101001";
                when "0000001001010" =>
                    dout1 <= "01101010";
                when "0000001001011" =>
                    dout1 <= "01101011";
                when "0000001001100" =>
                    dout1 <= "01101100";
                when "0000001001101" =>
                    dout1 <= "01101101";
                when "0000001001110" =>
                    dout1 <= "01101110";
                when "0000001001111" =>
                    dout1 <= "01101111";
                when "0000001010000" =>
                    dout1 <= "01110000";
                when "0000001010001" =>
                    dout1 <= "01110001";
                when "0000001010010" =>
                    dout1 <= "01110010";
                when "0000001010011" =>
                    dout1 <= "01110011";
                when "0000001010100" =>
                    dout1 <= "01110100";
                when "0000001010101" =>
                    dout1 <= "01110101";
                when "0000001010110" =>
                    dout1 <= "01110110";
                when "0000001010111" =>
                    dout1 <= "01110111";

    -- M global registers
                when "0000001011000" =>
                    dout1 <= "10000000";
                when "0000001011001" =>
                    dout1 <= "10000001";
                when "0000001011010" =>
                    dout1 <= "10000010";

        -- block #8

        -- 3*N registers for IN/LOC/OUT registers
                when "0000000100000" =>
                    dout1 <= "01110000";
                when "0000000100001" =>
                    dout1 <= "01110001";
                when "0000000100010" =>
                    dout1 <= "01110010";
                when "0000000100011" =>
                    dout1 <= "01110011";
                when "0000000100100" =>
                    dout1 <= "01110100";
                when "0000000100101" =>
                    dout1 <= "01110101";
                when "0000000100110" =>
                    dout1 <= "01110110";
                when "0000000100111" =>
                    dout1 <= "01110111";
                when "0000000101000" =>
                    dout1 <= "01111000";
                when "0000000101001" =>
                    dout1 <= "01111001";
                when "0000000101010" =>
                    dout1 <= "01111010";
                when "0000000101011" =>
                    dout1 <= "01111011";
                when "0000000101100" =>
                    dout1 <= "01111100";
                when "0000000101101" =>
                    dout1 <= "01111101";
                when "0000000101110" =>
                    dout1 <= "01111110";
                when "0000000101111" =>
                    dout1 <= "01111111";
                when "0000000110000" =>
                    dout1 <= "00000000";
                when "0000000110001" =>
                    dout1 <= "00000001";
                when "0000000110010" =>
                    dout1 <= "00000010";
                when "0000000110011" =>
                    dout1 <= "00000011";
                when "0000000110100" =>
                    dout1 <= "00000100";
                when "0000000110101" =>
                    dout1 <= "00000101";
                when "0000000110110" =>
                    dout1 <= "00000110";
                when "0000000110111" =>
                    dout1 <= "00000111";

    -- M global registers
                when "0000000111000" =>
                    dout1 <= "10000000";
                when "0000000111001" =>
                    dout1 <= "10000001";
                when "0000000111010" =>
                    dout1 <= "10000010";

    -- If enable not active the default output it 0
                when others =>
                    dout1 <= (others => '0');
            end case;
        end if;
    end process;

    -- Output port #2
    process(Clk, addr2, en)
        variable en_addr : std_logic_vector(8+5-1 downto 0);
    begin
        en_addr := en & addr2;
        if (rising_edge(Clk)) then 
            case (en_addr) is
        -- block #1

        -- 3*N registers for IN/LOC/OUT registers
                when "1000000000000" =>
                    dout2 <= "00000000";
                when "1000000000001" =>
                    dout2 <= "00000001";
                when "1000000000010" =>
                    dout2 <= "00000010";
                when "1000000000011" =>
                    dout2 <= "00000011";
                when "1000000000100" =>
                    dout2 <= "00000100";
                when "1000000000101" =>
                    dout2 <= "00000101";
                when "1000000000110" =>
                    dout2 <= "00000110";
                when "1000000000111" =>
                    dout2 <= "00000111";
                when "1000000001000" =>
                    dout2 <= "00001000";
                when "1000000001001" =>
                    dout2 <= "00001001";
                when "1000000001010" =>
                    dout2 <= "00001010";
                when "1000000001011" =>
                    dout2 <= "00001011";
                when "1000000001100" =>
                    dout2 <= "00001100";
                when "1000000001101" =>
                    dout2 <= "00001101";
                when "1000000001110" =>
                    dout2 <= "00001110";
                when "1000000001111" =>
                    dout2 <= "00001111";
                when "1000000010000" =>
                    dout2 <= "00010000";
                when "1000000010001" =>
                    dout2 <= "00010001";
                when "1000000010010" =>
                    dout2 <= "00010010";
                when "1000000010011" =>
                    dout2 <= "00010011";
                when "1000000010100" =>
                    dout2 <= "00010100";
                when "1000000010101" =>
                    dout2 <= "00010101";
                when "1000000010110" =>
                    dout2 <= "00010110";
                when "1000000010111" =>
                    dout2 <= "00010111";

    -- M global registers
                when "1000000011000" =>
                    dout2 <= "10000000";
                when "1000000011001" =>
                    dout2 <= "10000001";
                when "1000000011010" =>
                    dout2 <= "10000010";

        -- block #2

        -- 3*N registers for IN/LOC/OUT registers
                when "0100000000000" =>
                    dout2 <= "00010000";
                when "0100000000001" =>
                    dout2 <= "00010001";
                when "0100000000010" =>
                    dout2 <= "00010010";
                when "0100000000011" =>
                    dout2 <= "00010011";
                when "0100000000100" =>
                    dout2 <= "00010100";
                when "0100000000101" =>
                    dout2 <= "00010101";
                when "0100000000110" =>
                    dout2 <= "00010110";
                when "0100000000111" =>
                    dout2 <= "00010111";
                when "0100000001000" =>
                    dout2 <= "00011000";
                when "0100000001001" =>
                    dout2 <= "00011001";
                when "0100000001010" =>
                    dout2 <= "00011010";
                when "0100000001011" =>
                    dout2 <= "00011011";
                when "0100000001100" =>
                    dout2 <= "00011100";
                when "0100000001101" =>
                    dout2 <= "00011101";
                when "0100000001110" =>
                    dout2 <= "00011110";
                when "0100000001111" =>
                    dout2 <= "00011111";
                when "0100000010000" =>
                    dout2 <= "00100000";
                when "0100000010001" =>
                    dout2 <= "00100001";
                when "0100000010010" =>
                    dout2 <= "00100010";
                when "0100000010011" =>
                    dout2 <= "00100011";
                when "0100000010100" =>
                    dout2 <= "00100100";
                when "0100000010101" =>
                    dout2 <= "00100101";
                when "0100000010110" =>
                    dout2 <= "00100110";
                when "0100000010111" =>
                    dout2 <= "00100111";

    -- M global registers
                when "0100000011000" =>
                    dout2 <= "10000000";
                when "0100000011001" =>
                    dout2 <= "10000001";
                when "0100000011010" =>
                    dout2 <= "10000010";

        -- block #3

        -- 3*N registers for IN/LOC/OUT registers
                when "0010000000000" =>
                    dout2 <= "00100000";
                when "0010000000001" =>
                    dout2 <= "00100001";
                when "0010000000010" =>
                    dout2 <= "00100010";
                when "0010000000011" =>
                    dout2 <= "00100011";
                when "0010000000100" =>
                    dout2 <= "00100100";
                when "0010000000101" =>
                    dout2 <= "00100101";
                when "0010000000110" =>
                    dout2 <= "00100110";
                when "0010000000111" =>
                    dout2 <= "00100111";
                when "0010000001000" =>
                    dout2 <= "00101000";
                when "0010000001001" =>
                    dout2 <= "00101001";
                when "0010000001010" =>
                    dout2 <= "00101010";
                when "0010000001011" =>
                    dout2 <= "00101011";
                when "0010000001100" =>
                    dout2 <= "00101100";
                when "0010000001101" =>
                    dout2 <= "00101101";
                when "0010000001110" =>
                    dout2 <= "00101110";
                when "0010000001111" =>
                    dout2 <= "00101111";
                when "0010000010000" =>
                    dout2 <= "00110000";
                when "0010000010001" =>
                    dout2 <= "00110001";
                when "0010000010010" =>
                    dout2 <= "00110010";
                when "0010000010011" =>
                    dout2 <= "00110011";
                when "0010000010100" =>
                    dout2 <= "00110100";
                when "0010000010101" =>
                    dout2 <= "00110101";
                when "0010000010110" =>
                    dout2 <= "00110110";
                when "0010000010111" =>
                    dout2 <= "00110111";

    -- M global registers
                when "0010000011000" =>
                    dout2 <= "10000000";
                when "0010000011001" =>
                    dout2 <= "10000001";
                when "0010000011010" =>
                    dout2 <= "10000010";

        -- block #4

        -- 3*N registers for IN/LOC/OUT registers
                when "0001000000000" =>
                    dout2 <= "00110000";
                when "0001000000001" =>
                    dout2 <= "00110001";
                when "0001000000010" =>
                    dout2 <= "00110010";
                when "0001000000011" =>
                    dout2 <= "00110011";
                when "0001000000100" =>
                    dout2 <= "00110100";
                when "0001000000101" =>
                    dout2 <= "00110101";
                when "0001000000110" =>
                    dout2 <= "00110110";
                when "0001000000111" =>
                    dout2 <= "00110111";
                when "0001000001000" =>
                    dout2 <= "00111000";
                when "0001000001001" =>
                    dout2 <= "00111001";
                when "0001000001010" =>
                    dout2 <= "00111010";
                when "0001000001011" =>
                    dout2 <= "00111011";
                when "0001000001100" =>
                    dout2 <= "00111100";
                when "0001000001101" =>
                    dout2 <= "00111101";
                when "0001000001110" =>
                    dout2 <= "00111110";
                when "0001000001111" =>
                    dout2 <= "00111111";
                when "0001000010000" =>
                    dout2 <= "01000000";
                when "0001000010001" =>
                    dout2 <= "01000001";
                when "0001000010010" =>
                    dout2 <= "01000010";
                when "0001000010011" =>
                    dout2 <= "01000011";
                when "0001000010100" =>
                    dout2 <= "01000100";
                when "0001000010101" =>
                    dout2 <= "01000101";
                when "0001000010110" =>
                    dout2 <= "01000110";
                when "0001000010111" =>
                    dout2 <= "01000111";

    -- M global registers
                when "0001000011000" =>
                    dout2 <= "10000000";
                when "0001000011001" =>
                    dout2 <= "10000001";
                when "0001000011010" =>
                    dout2 <= "10000010";

        -- block #5

        -- 3*N registers for IN/LOC/OUT registers
                when "0000100000000" =>
                    dout2 <= "01000000";
                when "0000100000001" =>
                    dout2 <= "01000001";
                when "0000100000010" =>
                    dout2 <= "01000010";
                when "0000100000011" =>
                    dout2 <= "01000011";
                when "0000100000100" =>
                    dout2 <= "01000100";
                when "0000100000101" =>
                    dout2 <= "01000101";
                when "0000100000110" =>
                    dout2 <= "01000110";
                when "0000100000111" =>
                    dout2 <= "01000111";
                when "0000100001000" =>
                    dout2 <= "01001000";
                when "0000100001001" =>
                    dout2 <= "01001001";
                when "0000100001010" =>
                    dout2 <= "01001010";
                when "0000100001011" =>
                    dout2 <= "01001011";
                when "0000100001100" =>
                    dout2 <= "01001100";
                when "0000100001101" =>
                    dout2 <= "01001101";
                when "0000100001110" =>
                    dout2 <= "01001110";
                when "0000100001111" =>
                    dout2 <= "01001111";
                when "0000100010000" =>
                    dout2 <= "01010000";
                when "0000100010001" =>
                    dout2 <= "01010001";
                when "0000100010010" =>
                    dout2 <= "01010010";
                when "0000100010011" =>
                    dout2 <= "01010011";
                when "0000100010100" =>
                    dout2 <= "01010100";
                when "0000100010101" =>
                    dout2 <= "01010101";
                when "0000100010110" =>
                    dout2 <= "01010110";
                when "0000100010111" =>
                    dout2 <= "01010111";

    -- M global registers
                when "0000100011000" =>
                    dout2 <= "10000000";
                when "0000100011001" =>
                    dout2 <= "10000001";
                when "0000100011010" =>
                    dout2 <= "10000010";

        -- block #6

        -- 3*N registers for IN/LOC/OUT registers
                when "0000010000000" =>
                    dout2 <= "01010000";
                when "0000010000001" =>
                    dout2 <= "01010001";
                when "0000010000010" =>
                    dout2 <= "01010010";
                when "0000010000011" =>
                    dout2 <= "01010011";
                when "0000010000100" =>
                    dout2 <= "01010100";
                when "0000010000101" =>
                    dout2 <= "01010101";
                when "0000010000110" =>
                    dout2 <= "01010110";
                when "0000010000111" =>
                    dout2 <= "01010111";
                when "0000010001000" =>
                    dout2 <= "01011000";
                when "0000010001001" =>
                    dout2 <= "01011001";
                when "0000010001010" =>
                    dout2 <= "01011010";
                when "0000010001011" =>
                    dout2 <= "01011011";
                when "0000010001100" =>
                    dout2 <= "01011100";
                when "0000010001101" =>
                    dout2 <= "01011101";
                when "0000010001110" =>
                    dout2 <= "01011110";
                when "0000010001111" =>
                    dout2 <= "01011111";
                when "0000010010000" =>
                    dout2 <= "01100000";
                when "0000010010001" =>
                    dout2 <= "01100001";
                when "0000010010010" =>
                    dout2 <= "01100010";
                when "0000010010011" =>
                    dout2 <= "01100011";
                when "0000010010100" =>
                    dout2 <= "01100100";
                when "0000010010101" =>
                    dout2 <= "01100101";
                when "0000010010110" =>
                    dout2 <= "01100110";
                when "0000010010111" =>
                    dout2 <= "01100111";

    -- M global registers
                when "0000010011000" =>
                    dout2 <= "10000000";
                when "0000010011001" =>
                    dout2 <= "10000001";
                when "0000010011010" =>
                    dout2 <= "10000010";

        -- block #7

        -- 3*N registers for IN/LOC/OUT registers
                when "0000001000000" =>
                    dout2 <= "01100000";
                when "0000001000001" =>
                    dout2 <= "01100001";
                when "0000001000010" =>
                    dout2 <= "01100010";
                when "0000001000011" =>
                    dout2 <= "01100011";
                when "0000001000100" =>
                    dout2 <= "01100100";
                when "0000001000101" =>
                    dout2 <= "01100101";
                when "0000001000110" =>
                    dout2 <= "01100110";
                when "0000001000111" =>
                    dout2 <= "01100111";
                when "0000001001000" =>
                    dout2 <= "01101000";
                when "0000001001001" =>
                    dout2 <= "01101001";
                when "0000001001010" =>
                    dout2 <= "01101010";
                when "0000001001011" =>
                    dout2 <= "01101011";
                when "0000001001100" =>
                    dout2 <= "01101100";
                when "0000001001101" =>
                    dout2 <= "01101101";
                when "0000001001110" =>
                    dout2 <= "01101110";
                when "0000001001111" =>
                    dout2 <= "01101111";
                when "0000001010000" =>
                    dout2 <= "01110000";
                when "0000001010001" =>
                    dout2 <= "01110001";
                when "0000001010010" =>
                    dout2 <= "01110010";
                when "0000001010011" =>
                    dout2 <= "01110011";
                when "0000001010100" =>
                    dout2 <= "01110100";
                when "0000001010101" =>
                    dout2 <= "01110101";
                when "0000001010110" =>
                    dout2 <= "01110110";
                when "0000001010111" =>
                    dout2 <= "01110111";

    -- M global registers
                when "0000001011000" =>
                    dout2 <= "10000000";
                when "0000001011001" =>
                    dout2 <= "10000001";
                when "0000001011010" =>
                    dout2 <= "10000010";

        -- block #8

        -- 3*N registers for IN/LOC/OUT registers
                when "0000000100000" =>
                    dout2 <= "01110000";
                when "0000000100001" =>
                    dout2 <= "01110001";
                when "0000000100010" =>
                    dout2 <= "01110010";
                when "0000000100011" =>
                    dout2 <= "01110011";
                when "0000000100100" =>
                    dout2 <= "01110100";
                when "0000000100101" =>
                    dout2 <= "01110101";
                when "0000000100110" =>
                    dout2 <= "01110110";
                when "0000000100111" =>
                    dout2 <= "01110111";
                when "0000000101000" =>
                    dout2 <= "01111000";
                when "0000000101001" =>
                    dout2 <= "01111001";
                when "0000000101010" =>
                    dout2 <= "01111010";
                when "0000000101011" =>
                    dout2 <= "01111011";
                when "0000000101100" =>
                    dout2 <= "01111100";
                when "0000000101101" =>
                    dout2 <= "01111101";
                when "0000000101110" =>
                    dout2 <= "01111110";
                when "0000000101111" =>
                    dout2 <= "01111111";
                when "0000000110000" =>
                    dout2 <= "00000000";
                when "0000000110001" =>
                    dout2 <= "00000001";
                when "0000000110010" =>
                    dout2 <= "00000010";
                when "0000000110011" =>
                    dout2 <= "00000011";
                when "0000000110100" =>
                    dout2 <= "00000100";
                when "0000000110101" =>
                    dout2 <= "00000101";
                when "0000000110110" =>
                    dout2 <= "00000110";
                when "0000000110111" =>
                    dout2 <= "00000111";

    -- M global registers
                when "0000000111000" =>
                    dout2 <= "10000000";
                when "0000000111001" =>
                    dout2 <= "10000001";
                when "0000000111010" =>
                    dout2 <= "10000010";

    -- If enable not active the default output it 0
                when others =>
                    dout2 <= (others => '0');
            end case;
        end if;
    end process;
end architecture;

configuration CFG_LUT_ROM_ARCHBEH of LUT_ROM is
    for beh
    end for; 
end configuration;