
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_registerfile_M5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_registerfile_M5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerfile_M5.all;

entity registerfile_M5 is

   port( Clk, Rst, En, RD1, RD2, WR : in std_logic;  Addr_WR, Addr_RD1, 
         Addr_RD2 : in std_logic_vector (4 downto 0);  DataIN : in 
         std_logic_vector (31 downto 0);  Out1, Out2 : out std_logic_vector (31
         downto 0));

end registerfile_M5;

architecture SYN_ARCHBEH of registerfile_M5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal Out1_31_port, Out1_30_port, Out1_29_port, Out1_28_port, Out1_27_port,
      Out1_26_port, Out1_25_port, Out1_24_port, Out1_23_port, Out1_22_port, 
      Out1_21_port, Out1_20_port, Out1_19_port, Out1_18_port, Out1_17_port, 
      Out1_16_port, Out1_15_port, Out1_14_port, Out1_13_port, Out1_12_port, 
      Out1_11_port, Out1_10_port, Out1_9_port, Out1_8_port, Out1_7_port, 
      Out1_6_port, Out1_5_port, Out1_4_port, Out1_3_port, Out1_2_port, 
      Out1_1_port, Out1_0_port, Out2_31_port, Out2_30_port, Out2_29_port, 
      Out2_28_port, Out2_27_port, Out2_26_port, Out2_25_port, Out2_24_port, 
      Out2_23_port, Out2_22_port, Out2_21_port, Out2_20_port, Out2_19_port, 
      Out2_18_port, Out2_17_port, Out2_16_port, Out2_15_port, Out2_14_port, 
      Out2_13_port, Out2_12_port, Out2_11_port, Out2_10_port, Out2_9_port, 
      Out2_8_port, Out2_7_port, Out2_6_port, Out2_5_port, Out2_4_port, 
      Out2_3_port, Out2_2_port, Out2_1_port, Out2_0_port, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, 
      n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, 
      n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
      n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
      n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
      n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, 
      n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
      n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
      n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
      n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
      n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
      n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, 
      n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, 
      n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, 
      n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, 
      n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, 
      n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, 
      n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, 
      n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
      n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, 
      n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
      n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, 
      n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, 
      n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, 
      n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, 
      n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
      n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, 
      n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, 
      n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
      n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
      n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
      n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, 
      n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, 
      n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, 
      n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, 
      n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, 
      n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, 
      n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, 
      n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
      n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, 
      n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
      n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, 
      n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
      n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, 
      n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
      n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
      n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
      n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, 
      n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
      n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
      n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
      n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
      n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
      n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
      n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
      n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
      n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, 
      n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
      n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
      n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, 
      n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, 
      n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
      n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
      n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, 
      n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
      n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
      n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, 
      n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, 
      n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, 
      n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, 
      n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, 
      n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, 
      n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, 
      n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, 
      n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
      n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, 
      n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, 
      n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, 
      n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
      n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, 
      n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
      n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
      n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
      n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
      n2301, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, 
      n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, 
      n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, 
      n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, 
      n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, 
      n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, 
      n7273, n7274, n7275, n7276, n7277, n7374, n7375, n7376, n7377, n7378, 
      n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, 
      n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, 
      n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7470, n7471, n7472, 
      n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, 
      n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, 
      n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7534, 
      n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, 
      n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, 
      n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, 
      n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, 
      n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, 
      n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, 
      n7595, n7596, n7597, n8260, n8261, n8262, n8263, n8264, n8265, n8266, 
      n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, 
      n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, 
      n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, 
      n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, 
      n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, 
      n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, 
      n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, 
      n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, 
      n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, 
      n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, 
      n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, 
      n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, 
      n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, 
      n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, 
      n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, 
      n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, 
      n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, 
      n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, 
      n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, 
      n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, 
      n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, 
      n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, 
      n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, 
      n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, 
      n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, 
      n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, 
      n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, 
      n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, 
      n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, 
      n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, 
      n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, 
      n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, 
      n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, 
      n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, 
      n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, 
      n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, 
      n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, 
      n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, 
      n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, 
      n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, 
      n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, 
      n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, 
      n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, 
      n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, 
      n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, 
      n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, 
      n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, 
      n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, 
      n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, 
      n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, 
      n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, 
      n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, 
      n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, 
      n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, 
      n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, 
      n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, 
      n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, 
      n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, 
      n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, 
      n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, 
      n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, 
      n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, 
      n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, 
      n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, 
      n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, 
      n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, 
      n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, 
      n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, 
      n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, 
      n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, 
      n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, 
      n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, 
      n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, 
      n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, 
      n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, 
      n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, 
      n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, 
      n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, 
      n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, 
      n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, 
      n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, 
      n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, 
      n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, 
      n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, 
      n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, 
      n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, 
      n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, 
      n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, 
      n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, 
      n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, 
      n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, 
      n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, 
      n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, 
      n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, 
      n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, 
      n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, 
      n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, 
      n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, 
      n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, 
      n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, 
      n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, 
      n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, 
      n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, 
      n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, 
      n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, 
      n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, 
      n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, 
      n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, 
      n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, 
      n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, 
      n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, 
      n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, 
      n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, 
      n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, 
      n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, 
      n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, 
      n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, 
      n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, 
      n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, 
      n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, 
      n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, 
      n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, 
      n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, 
      n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, 
      n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, 
      n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, 
      n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, 
      n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, 
      n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, 
      n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, 
      n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, 
      n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, 
      n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, 
      n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, 
      n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, 
      n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, 
      n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, 
      n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, 
      n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, 
      n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, 
      n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, 
      n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, 
      n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, 
      n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, 
      n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, 
      n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, 
      n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, 
      n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, 
      n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, 
      n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, 
      n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, 
      n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, 
      n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, 
      n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, 
      n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, 
      n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, 
      n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, 
      n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, 
      n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, 
      n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, 
      n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, 
      n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, 
      n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, 
      n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, 
      n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, 
      n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, 
      n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, 
      n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, 
      n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, 
      n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, 
      n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, 
      n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, 
      n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, 
      n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, 
      n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, 
      n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, 
      n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, 
      n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, 
      n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, 
      n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, 
      n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, 
      n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, 
      n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, 
      n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, 
      n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, 
      n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, 
      n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, 
      n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, 
      n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, 
      n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, 
      n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, 
      n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, 
      n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, 
      n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, 
      n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, 
      n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, 
      n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, 
      n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, 
      n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, 
      n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, 
      n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, 
      n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, 
      n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, 
      n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, 
      n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, 
      n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, 
      n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, 
      n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, 
      n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, 
      n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, 
      n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, 
      n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, 
      n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, 
      n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, 
      n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, 
      n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, 
      n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, 
      n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, 
      n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, 
      n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, 
      n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, 
      n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, 
      n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, 
      n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, 
      n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, 
      n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, 
      n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, 
      n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, 
      n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, 
      n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, 
      n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, 
      n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, 
      n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, 
      n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, 
      n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, 
      n10555, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, 
      n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, 
      n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, 
      n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, 
      n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, 
      n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, 
      n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, 
      n10747, n10748, n10845, n10846, n10847, n10848, n10849, n10850, n10851, 
      n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, 
      n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, 
      n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10909, n10910, 
      n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, 
      n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, 
      n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, 
      n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, 
      n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, 
      n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, 
      n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, 
      n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, 
      n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, 
      n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, 
      n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, 
      n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, 
      n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, 
      n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, 
      n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, 
      n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, 
      n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, 
      n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, 
      n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, 
      n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, 
      n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, 
      n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, 
      n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, 
      n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, 
      n11191, n11192, n11193, n11194, n11195, n11196, n11260, n11261, n11262, 
      n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, 
      n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, 
      n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, 
      n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, 
      n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, 
      n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, 
      n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, 
      n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, 
      n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, 
      n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, 
      n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, 
      n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, 
      n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, 
      n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, 
      n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, 
      n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, 
      n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, 
      n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, 
      n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, 
      n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, 
      n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, 
      n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, 
      n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, 
      n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, 
      n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, 
      n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, 
      n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, 
      n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, 
      n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, 
      n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, 
      n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, 
      n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, 
      n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, 
      n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, 
      n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, 
      n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, 
      n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, 
      n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, 
      n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, 
      n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, 
      n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, 
      n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, 
      n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, 
      n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, 
      n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, 
      n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, 
      n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, 
      n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, 
      n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, 
      n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, 
      n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, 
      n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, 
      n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, 
      n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, 
      n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, 
      n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, 
      n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, 
      n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, 
      n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, 
      n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, 
      n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, 
      n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, 
      n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, 
      n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, 
      n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, 
      n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, 
      n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, 
      n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, 
      n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, 
      n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, 
      n11893, n11894, n11895, n11896, n11897, n_1000, n_1001, n_1002, n_1003, 
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639 : std_logic;

begin
   Out1 <= ( Out1_31_port, Out1_30_port, Out1_29_port, Out1_28_port, 
      Out1_27_port, Out1_26_port, Out1_25_port, Out1_24_port, Out1_23_port, 
      Out1_22_port, Out1_21_port, Out1_20_port, Out1_19_port, Out1_18_port, 
      Out1_17_port, Out1_16_port, Out1_15_port, Out1_14_port, Out1_13_port, 
      Out1_12_port, Out1_11_port, Out1_10_port, Out1_9_port, Out1_8_port, 
      Out1_7_port, Out1_6_port, Out1_5_port, Out1_4_port, Out1_3_port, 
      Out1_2_port, Out1_1_port, Out1_0_port );
   Out2 <= ( Out2_31_port, Out2_30_port, Out2_29_port, Out2_28_port, 
      Out2_27_port, Out2_26_port, Out2_25_port, Out2_24_port, Out2_23_port, 
      Out2_22_port, Out2_21_port, Out2_20_port, Out2_19_port, Out2_18_port, 
      Out2_17_port, Out2_16_port, Out2_15_port, Out2_14_port, Out2_13_port, 
      Out2_12_port, Out2_11_port, Out2_10_port, Out2_9_port, Out2_8_port, 
      Out2_7_port, Out2_6_port, Out2_5_port, Out2_4_port, Out2_3_port, 
      Out2_2_port, Out2_1_port, Out2_0_port );
   
   Out1_reg_31_inst : DFF_X1 port map( D => n7277, CK => Clk, Q => Out1_31_port
                           , QN => n_1000);
   Out1_reg_30_inst : DFF_X1 port map( D => n7276, CK => Clk, Q => Out1_30_port
                           , QN => n_1001);
   Out1_reg_29_inst : DFF_X1 port map( D => n7275, CK => Clk, Q => Out1_29_port
                           , QN => n_1002);
   Out1_reg_28_inst : DFF_X1 port map( D => n7274, CK => Clk, Q => Out1_28_port
                           , QN => n_1003);
   Out1_reg_27_inst : DFF_X1 port map( D => n7273, CK => Clk, Q => Out1_27_port
                           , QN => n_1004);
   Out1_reg_26_inst : DFF_X1 port map( D => n7272, CK => Clk, Q => Out1_26_port
                           , QN => n_1005);
   Out1_reg_25_inst : DFF_X1 port map( D => n7271, CK => Clk, Q => Out1_25_port
                           , QN => n_1006);
   Out1_reg_24_inst : DFF_X1 port map( D => n7270, CK => Clk, Q => Out1_24_port
                           , QN => n_1007);
   Out1_reg_23_inst : DFF_X1 port map( D => n7269, CK => Clk, Q => Out1_23_port
                           , QN => n_1008);
   Out1_reg_22_inst : DFF_X1 port map( D => n7268, CK => Clk, Q => Out1_22_port
                           , QN => n_1009);
   Out1_reg_21_inst : DFF_X1 port map( D => n7267, CK => Clk, Q => Out1_21_port
                           , QN => n_1010);
   Out1_reg_20_inst : DFF_X1 port map( D => n7266, CK => Clk, Q => Out1_20_port
                           , QN => n_1011);
   Out1_reg_19_inst : DFF_X1 port map( D => n7265, CK => Clk, Q => Out1_19_port
                           , QN => n_1012);
   Out1_reg_18_inst : DFF_X1 port map( D => n7264, CK => Clk, Q => Out1_18_port
                           , QN => n_1013);
   Out1_reg_17_inst : DFF_X1 port map( D => n7263, CK => Clk, Q => Out1_17_port
                           , QN => n_1014);
   Out1_reg_16_inst : DFF_X1 port map( D => n7262, CK => Clk, Q => Out1_16_port
                           , QN => n_1015);
   Out1_reg_15_inst : DFF_X1 port map( D => n7261, CK => Clk, Q => Out1_15_port
                           , QN => n_1016);
   Out1_reg_14_inst : DFF_X1 port map( D => n7260, CK => Clk, Q => Out1_14_port
                           , QN => n_1017);
   Out1_reg_13_inst : DFF_X1 port map( D => n7259, CK => Clk, Q => Out1_13_port
                           , QN => n_1018);
   Out1_reg_12_inst : DFF_X1 port map( D => n7258, CK => Clk, Q => Out1_12_port
                           , QN => n_1019);
   Out1_reg_11_inst : DFF_X1 port map( D => n7257, CK => Clk, Q => Out1_11_port
                           , QN => n_1020);
   Out1_reg_10_inst : DFF_X1 port map( D => n7256, CK => Clk, Q => Out1_10_port
                           , QN => n_1021);
   Out1_reg_9_inst : DFF_X1 port map( D => n7255, CK => Clk, Q => Out1_9_port, 
                           QN => n_1022);
   Out1_reg_8_inst : DFF_X1 port map( D => n7254, CK => Clk, Q => Out1_8_port, 
                           QN => n_1023);
   Out1_reg_7_inst : DFF_X1 port map( D => n7253, CK => Clk, Q => Out1_7_port, 
                           QN => n_1024);
   Out1_reg_6_inst : DFF_X1 port map( D => n7252, CK => Clk, Q => Out1_6_port, 
                           QN => n_1025);
   Out1_reg_5_inst : DFF_X1 port map( D => n7251, CK => Clk, Q => Out1_5_port, 
                           QN => n_1026);
   Out1_reg_4_inst : DFF_X1 port map( D => n7250, CK => Clk, Q => Out1_4_port, 
                           QN => n_1027);
   Out1_reg_3_inst : DFF_X1 port map( D => n7249, CK => Clk, Q => Out1_3_port, 
                           QN => n_1028);
   Out1_reg_2_inst : DFF_X1 port map( D => n7248, CK => Clk, Q => Out1_2_port, 
                           QN => n_1029);
   Out1_reg_1_inst : DFF_X1 port map( D => n7247, CK => Clk, Q => Out1_1_port, 
                           QN => n_1030);
   Out1_reg_0_inst : DFF_X1 port map( D => n7246, CK => Clk, Q => Out1_0_port, 
                           QN => n_1031);
   Out2_reg_30_inst : DFF_X1 port map( D => n7244, CK => Clk, Q => Out2_30_port
                           , QN => n_1032);
   Out2_reg_29_inst : DFF_X1 port map( D => n7243, CK => Clk, Q => Out2_29_port
                           , QN => n_1033);
   Out2_reg_28_inst : DFF_X1 port map( D => n7242, CK => Clk, Q => Out2_28_port
                           , QN => n_1034);
   Out2_reg_27_inst : DFF_X1 port map( D => n7241, CK => Clk, Q => Out2_27_port
                           , QN => n_1035);
   Out2_reg_26_inst : DFF_X1 port map( D => n7240, CK => Clk, Q => Out2_26_port
                           , QN => n_1036);
   Out2_reg_25_inst : DFF_X1 port map( D => n7239, CK => Clk, Q => Out2_25_port
                           , QN => n_1037);
   Out2_reg_24_inst : DFF_X1 port map( D => n7238, CK => Clk, Q => Out2_24_port
                           , QN => n_1038);
   Out2_reg_23_inst : DFF_X1 port map( D => n7237, CK => Clk, Q => Out2_23_port
                           , QN => n_1039);
   Out2_reg_22_inst : DFF_X1 port map( D => n7236, CK => Clk, Q => Out2_22_port
                           , QN => n_1040);
   Out2_reg_21_inst : DFF_X1 port map( D => n7235, CK => Clk, Q => Out2_21_port
                           , QN => n_1041);
   Out2_reg_20_inst : DFF_X1 port map( D => n7234, CK => Clk, Q => Out2_20_port
                           , QN => n_1042);
   Out2_reg_19_inst : DFF_X1 port map( D => n7233, CK => Clk, Q => Out2_19_port
                           , QN => n_1043);
   Out2_reg_18_inst : DFF_X1 port map( D => n7232, CK => Clk, Q => Out2_18_port
                           , QN => n_1044);
   Out2_reg_17_inst : DFF_X1 port map( D => n7231, CK => Clk, Q => Out2_17_port
                           , QN => n_1045);
   Out2_reg_16_inst : DFF_X1 port map( D => n7230, CK => Clk, Q => Out2_16_port
                           , QN => n_1046);
   Out2_reg_15_inst : DFF_X1 port map( D => n7229, CK => Clk, Q => Out2_15_port
                           , QN => n_1047);
   Out2_reg_14_inst : DFF_X1 port map( D => n7228, CK => Clk, Q => Out2_14_port
                           , QN => n_1048);
   Out2_reg_13_inst : DFF_X1 port map( D => n7227, CK => Clk, Q => Out2_13_port
                           , QN => n_1049);
   Out2_reg_12_inst : DFF_X1 port map( D => n7226, CK => Clk, Q => Out2_12_port
                           , QN => n_1050);
   Out2_reg_11_inst : DFF_X1 port map( D => n7225, CK => Clk, Q => Out2_11_port
                           , QN => n_1051);
   Out2_reg_10_inst : DFF_X1 port map( D => n7224, CK => Clk, Q => Out2_10_port
                           , QN => n_1052);
   Out2_reg_9_inst : DFF_X1 port map( D => n7223, CK => Clk, Q => Out2_9_port, 
                           QN => n_1053);
   Out2_reg_8_inst : DFF_X1 port map( D => n7222, CK => Clk, Q => Out2_8_port, 
                           QN => n_1054);
   Out2_reg_7_inst : DFF_X1 port map( D => n7221, CK => Clk, Q => Out2_7_port, 
                           QN => n_1055);
   Out2_reg_6_inst : DFF_X1 port map( D => n7220, CK => Clk, Q => Out2_6_port, 
                           QN => n_1056);
   Out2_reg_5_inst : DFF_X1 port map( D => n7219, CK => Clk, Q => Out2_5_port, 
                           QN => n_1057);
   Out2_reg_4_inst : DFF_X1 port map( D => n7218, CK => Clk, Q => Out2_4_port, 
                           QN => n_1058);
   Out2_reg_3_inst : DFF_X1 port map( D => n7217, CK => Clk, Q => Out2_3_port, 
                           QN => n_1059);
   Out2_reg_2_inst : DFF_X1 port map( D => n7216, CK => Clk, Q => Out2_2_port, 
                           QN => n_1060);
   Out2_reg_1_inst : DFF_X1 port map( D => n7215, CK => Clk, Q => Out2_1_port, 
                           QN => n_1061);
   Out2_reg_0_inst : DFF_X1 port map( D => n7214, CK => Clk, Q => Out2_0_port, 
                           QN => n_1062);
   U7498 : NAND3_X1 port map( A1 => n9864, A2 => n11838, A3 => n9865, ZN => 
                           n9306);
   U7499 : NAND3_X1 port map( A1 => n9866, A2 => n11838, A3 => n9867, ZN => 
                           n9305);
   U7500 : NAND3_X1 port map( A1 => n9865, A2 => n11838, A3 => n9868, ZN => 
                           n9311);
   U7501 : NAND3_X1 port map( A1 => n9865, A2 => n11838, A3 => n9870, ZN => 
                           n9310);
   U7502 : NAND3_X1 port map( A1 => n9867, A2 => n11838, A3 => n9870, ZN => 
                           n9316);
   U7503 : NAND3_X1 port map( A1 => n9867, A2 => n11838, A3 => n9873, ZN => 
                           n9315);
   U7504 : NAND3_X1 port map( A1 => n9865, A2 => n11838, A3 => n9871, ZN => 
                           n9322);
   U7505 : NAND3_X1 port map( A1 => n9867, A2 => n11838, A3 => n9874, ZN => 
                           n9321);
   U7506 : NAND3_X1 port map( A1 => n10454, A2 => n11699, A3 => n10455, ZN => 
                           n9896);
   U7507 : NAND3_X1 port map( A1 => n10456, A2 => n11699, A3 => n10457, ZN => 
                           n9895);
   U7508 : NAND3_X1 port map( A1 => n10455, A2 => n11699, A3 => n10458, ZN => 
                           n9901);
   U7509 : NAND3_X1 port map( A1 => n10455, A2 => n11699, A3 => n10460, ZN => 
                           n9900);
   U7510 : NAND3_X1 port map( A1 => n10457, A2 => n11699, A3 => n10460, ZN => 
                           n9906);
   U7511 : NAND3_X1 port map( A1 => n10457, A2 => n11699, A3 => n10463, ZN => 
                           n9905);
   U7512 : NAND3_X1 port map( A1 => n10455, A2 => n11699, A3 => n10461, ZN => 
                           n9912);
   U7513 : NAND3_X1 port map( A1 => n10457, A2 => n11699, A3 => n10464, ZN => 
                           n9911);
   U7514 : NAND3_X1 port map( A1 => n8263, A2 => n8262, A3 => n10519, ZN => 
                           n10511);
   U7515 : NAND3_X1 port map( A1 => n10519, A2 => n8262, A3 => Addr_WR(2), ZN 
                           => n10521);
   U7516 : NAND3_X1 port map( A1 => n10519, A2 => n8263, A3 => Addr_WR(3), ZN 
                           => n10526);
   U7517 : NAND3_X1 port map( A1 => Addr_WR(2), A2 => n10519, A3 => Addr_WR(3),
                           ZN => n10531);
   U7518 : NAND3_X1 port map( A1 => n8263, A2 => n8262, A3 => n10540, ZN => 
                           n10536);
   U7519 : NAND3_X1 port map( A1 => Addr_WR(2), A2 => n8262, A3 => n10540, ZN 
                           => n10542);
   U7520 : NAND3_X1 port map( A1 => Addr_WR(3), A2 => n8263, A3 => n10540, ZN 
                           => n10547);
   U7521 : NAND3_X1 port map( A1 => Addr_WR(3), A2 => Addr_WR(2), A3 => n10540,
                           ZN => n10552);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1309, CK => Clk, Q => 
                           n_1063, QN => n9266);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1308, CK => Clk, Q => 
                           n_1064, QN => n9267);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1307, CK => Clk, Q => 
                           n_1065, QN => n9268);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1306, CK => Clk, Q => 
                           n_1066, QN => n9269);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1305, CK => Clk, Q => 
                           n_1067, QN => n9270);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1304, CK => Clk, Q => 
                           n_1068, QN => n9271);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1303, CK => Clk, Q => 
                           n_1069, QN => n9272);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1302, CK => Clk, Q => 
                           n_1070, QN => n9273);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1301, CK => Clk, Q => 
                           n_1071, QN => n9274);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1300, CK => Clk, Q => 
                           n_1072, QN => n9275);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1299, CK => Clk, Q => 
                           n_1073, QN => n9276);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1298, CK => Clk, Q => 
                           n_1074, QN => n9277);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1297, CK => Clk, Q => 
                           n_1075, QN => n9278);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1296, CK => Clk, Q => 
                           n_1076, QN => n9279);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1295, CK => Clk, Q => 
                           n_1077, QN => n9280);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1294, CK => Clk, Q => 
                           n_1078, QN => n9281);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1293, CK => Clk, Q => 
                           n_1079, QN => n9282);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1292, CK => Clk, Q => 
                           n_1080, QN => n9283);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1291, CK => Clk, Q => 
                           n_1081, QN => n9284);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1290, CK => Clk, Q => 
                           n_1082, QN => n9285);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1289, CK => Clk, Q => 
                           n_1083, QN => n9286);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1288, CK => Clk, Q => 
                           n_1084, QN => n9287);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1287, CK => Clk, Q => 
                           n_1085, QN => n9288);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1286, CK => Clk, Q => 
                           n_1086, QN => n9289);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1285, CK => Clk, Q => 
                           n_1087, QN => n9290);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1284, CK => Clk, Q => 
                           n_1088, QN => n9291);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1283, CK => Clk, Q => 
                           n_1089, QN => n9292);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1282, CK => Clk, Q => 
                           n_1090, QN => n9293);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1281, CK => Clk, Q => 
                           n_1091, QN => n9294);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1280, CK => Clk, Q => 
                           n_1092, QN => n9295);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1279, CK => Clk, Q => 
                           n_1093, QN => n9296);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1278, CK => Clk, Q => 
                           n_1094, QN => n9297);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1981, CK => Clk, Q => 
                           n_1095, QN => n8594);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1980, CK => Clk, Q => 
                           n_1096, QN => n8595);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1979, CK => Clk, Q => 
                           n_1097, QN => n8596);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1978, CK => Clk, Q => 
                           n_1098, QN => n8597);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1977, CK => Clk, Q => 
                           n_1099, QN => n8598);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1976, CK => Clk, Q => 
                           n_1100, QN => n8599);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1975, CK => Clk, Q => 
                           n_1101, QN => n8600);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1974, CK => Clk, Q => 
                           n_1102, QN => n8601);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2269, CK => Clk, Q => 
                           n_1103, QN => n8306);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2268, CK => Clk, Q => 
                           n_1104, QN => n8307);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2267, CK => Clk, Q => 
                           n_1105, QN => n8308);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2266, CK => Clk, Q => 
                           n_1106, QN => n8309);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2265, CK => Clk, Q => 
                           n_1107, QN => n8310);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2264, CK => Clk, Q => 
                           n_1108, QN => n8311);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2263, CK => Clk, Q => 
                           n_1109, QN => n8312);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2262, CK => Clk, Q => 
                           n_1110, QN => n8313);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1973, CK => Clk, Q => 
                           n_1111, QN => n8602);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1972, CK => Clk, Q => 
                           n_1112, QN => n8603);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1971, CK => Clk, Q => 
                           n_1113, QN => n8604);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1970, CK => Clk, Q => 
                           n_1114, QN => n8605);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1969, CK => Clk, Q => 
                           n_1115, QN => n8606);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1968, CK => Clk, Q => 
                           n_1116, QN => n8607);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1967, CK => Clk, Q => 
                           n_1117, QN => n8608);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1966, CK => Clk, Q => 
                           n_1118, QN => n8609);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1965, CK => Clk, Q => 
                           n_1119, QN => n8610);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1964, CK => Clk, Q => 
                           n_1120, QN => n8611);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1963, CK => Clk, Q => 
                           n_1121, QN => n8612);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1962, CK => Clk, Q => 
                           n_1122, QN => n8613);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1961, CK => Clk, Q => 
                           n_1123, QN => n8614);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1960, CK => Clk, Q => 
                           n_1124, QN => n8615);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1959, CK => Clk, Q => 
                           n_1125, QN => n8616);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1958, CK => Clk, Q => 
                           n_1126, QN => n8617);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1957, CK => Clk, Q => 
                           n_1127, QN => n8618);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1956, CK => Clk, Q => 
                           n_1128, QN => n8619);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1955, CK => Clk, Q => 
                           n_1129, QN => n8620);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1954, CK => Clk, Q => 
                           n_1130, QN => n8621);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1953, CK => Clk, Q => 
                           n_1131, QN => n8622);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1952, CK => Clk, Q => 
                           n_1132, QN => n8623);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1951, CK => Clk, Q => 
                           n_1133, QN => n8624);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1950, CK => Clk, Q => 
                           n_1134, QN => n8625);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2261, CK => Clk, Q => 
                           n_1135, QN => n8314);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2260, CK => Clk, Q => 
                           n_1136, QN => n8315);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2259, CK => Clk, Q => 
                           n_1137, QN => n8316);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2258, CK => Clk, Q => 
                           n_1138, QN => n8317);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2257, CK => Clk, Q => 
                           n_1139, QN => n8318);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2256, CK => Clk, Q => 
                           n_1140, QN => n8319);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2255, CK => Clk, Q => 
                           n_1141, QN => n8320);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2254, CK => Clk, Q => 
                           n_1142, QN => n8321);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2253, CK => Clk, Q => 
                           n_1143, QN => n8322);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2252, CK => Clk, Q => 
                           n_1144, QN => n8323);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2251, CK => Clk, Q => 
                           n_1145, QN => n8324);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2250, CK => Clk, Q => 
                           n_1146, QN => n8325);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2249, CK => Clk, Q => 
                           n_1147, QN => n8326);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2248, CK => Clk, Q => 
                           n_1148, QN => n8327);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2247, CK => Clk, Q => n_1149
                           , QN => n8328);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2246, CK => Clk, Q => n_1150
                           , QN => n8329);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2245, CK => Clk, Q => n_1151
                           , QN => n8330);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2244, CK => Clk, Q => n_1152
                           , QN => n8331);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2243, CK => Clk, Q => n_1153
                           , QN => n8332);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2242, CK => Clk, Q => n_1154
                           , QN => n8333);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2241, CK => Clk, Q => n_1155
                           , QN => n8334);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2240, CK => Clk, Q => n_1156
                           , QN => n8335);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2239, CK => Clk, Q => n_1157
                           , QN => n8336);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2238, CK => Clk, Q => n_1158
                           , QN => n8337);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1341, CK => Clk, Q => 
                           n_1159, QN => n9234);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1340, CK => Clk, Q => 
                           n_1160, QN => n9235);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1339, CK => Clk, Q => 
                           n_1161, QN => n9236);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1338, CK => Clk, Q => 
                           n_1162, QN => n9237);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1337, CK => Clk, Q => 
                           n_1163, QN => n9238);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1336, CK => Clk, Q => 
                           n_1164, QN => n9239);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1335, CK => Clk, Q => 
                           n_1165, QN => n9240);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1334, CK => Clk, Q => 
                           n_1166, QN => n9241);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1501, CK => Clk, Q => 
                           n_1167, QN => n9074);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1500, CK => Clk, Q => 
                           n_1168, QN => n9075);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1499, CK => Clk, Q => 
                           n_1169, QN => n9076);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1498, CK => Clk, Q => 
                           n_1170, QN => n9077);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1497, CK => Clk, Q => 
                           n_1171, QN => n9078);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1496, CK => Clk, Q => 
                           n_1172, QN => n9079);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1495, CK => Clk, Q => 
                           n_1173, QN => n9080);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1494, CK => Clk, Q => 
                           n_1174, QN => n9081);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1629, CK => Clk, Q => 
                           n_1175, QN => n8946);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1628, CK => Clk, Q => 
                           n_1176, QN => n8947);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1627, CK => Clk, Q => 
                           n_1177, QN => n8948);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1626, CK => Clk, Q => 
                           n_1178, QN => n8949);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1625, CK => Clk, Q => 
                           n_1179, QN => n8950);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1624, CK => Clk, Q => 
                           n_1180, QN => n8951);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1623, CK => Clk, Q => 
                           n_1181, QN => n8952);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1622, CK => Clk, Q => 
                           n_1182, QN => n8953);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1661, CK => Clk, Q => 
                           n_1183, QN => n8914);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1660, CK => Clk, Q => 
                           n_1184, QN => n8915);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1659, CK => Clk, Q => 
                           n_1185, QN => n8916);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1658, CK => Clk, Q => 
                           n_1186, QN => n8917);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1657, CK => Clk, Q => 
                           n_1187, QN => n8918);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1656, CK => Clk, Q => 
                           n_1188, QN => n8919);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1655, CK => Clk, Q => 
                           n_1189, QN => n8920);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1654, CK => Clk, Q => 
                           n_1190, QN => n8921);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1949, CK => Clk, Q => 
                           n_1191, QN => n8626);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1948, CK => Clk, Q => 
                           n_1192, QN => n8627);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1947, CK => Clk, Q => 
                           n_1193, QN => n8628);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1946, CK => Clk, Q => 
                           n_1194, QN => n8629);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1945, CK => Clk, Q => 
                           n_1195, QN => n8630);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1944, CK => Clk, Q => 
                           n_1196, QN => n8631);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1943, CK => Clk, Q => 
                           n_1197, QN => n8632);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1942, CK => Clk, Q => 
                           n_1198, QN => n8633);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1885, CK => Clk, Q => 
                           n_1199, QN => n8690);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1884, CK => Clk, Q => 
                           n_1200, QN => n8691);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1883, CK => Clk, Q => 
                           n_1201, QN => n8692);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1882, CK => Clk, Q => 
                           n_1202, QN => n8693);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1881, CK => Clk, Q => 
                           n_1203, QN => n8694);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1880, CK => Clk, Q => 
                           n_1204, QN => n8695);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1879, CK => Clk, Q => 
                           n_1205, QN => n8696);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1878, CK => Clk, Q => 
                           n_1206, QN => n8697);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2237, CK => Clk, Q => 
                           n_1207, QN => n8338);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2236, CK => Clk, Q => 
                           n_1208, QN => n8339);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2235, CK => Clk, Q => 
                           n_1209, QN => n8340);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2234, CK => Clk, Q => 
                           n_1210, QN => n8341);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2233, CK => Clk, Q => 
                           n_1211, QN => n8342);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2232, CK => Clk, Q => 
                           n_1212, QN => n8343);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2231, CK => Clk, Q => 
                           n_1213, QN => n8344);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2230, CK => Clk, Q => 
                           n_1214, QN => n8345);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1373, CK => Clk, Q => 
                           n_1215, QN => n9202);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1372, CK => Clk, Q => 
                           n_1216, QN => n9203);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1371, CK => Clk, Q => 
                           n_1217, QN => n9204);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1370, CK => Clk, Q => 
                           n_1218, QN => n9205);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1369, CK => Clk, Q => 
                           n_1219, QN => n9206);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1368, CK => Clk, Q => 
                           n_1220, QN => n9207);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1367, CK => Clk, Q => 
                           n_1221, QN => n9208);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1366, CK => Clk, Q => 
                           n_1222, QN => n9209);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1405, CK => Clk, Q => 
                           n_1223, QN => n9170);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1404, CK => Clk, Q => 
                           n_1224, QN => n9171);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1403, CK => Clk, Q => 
                           n_1225, QN => n9172);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1402, CK => Clk, Q => 
                           n_1226, QN => n9173);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1401, CK => Clk, Q => 
                           n_1227, QN => n9174);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1400, CK => Clk, Q => 
                           n_1228, QN => n9175);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1399, CK => Clk, Q => 
                           n_1229, QN => n9176);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1398, CK => Clk, Q => 
                           n_1230, QN => n9177);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1693, CK => Clk, Q => 
                           n_1231, QN => n8882);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1692, CK => Clk, Q => 
                           n_1232, QN => n8883);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1691, CK => Clk, Q => 
                           n_1233, QN => n8884);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1690, CK => Clk, Q => 
                           n_1234, QN => n8885);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1689, CK => Clk, Q => 
                           n_1235, QN => n8886);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1688, CK => Clk, Q => 
                           n_1236, QN => n8887);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1687, CK => Clk, Q => 
                           n_1237, QN => n8888);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1686, CK => Clk, Q => 
                           n_1238, QN => n8889);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1725, CK => Clk, Q => 
                           n_1239, QN => n8850);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1724, CK => Clk, Q => 
                           n_1240, QN => n8851);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1723, CK => Clk, Q => 
                           n_1241, QN => n8852);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1722, CK => Clk, Q => 
                           n_1242, QN => n8853);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1721, CK => Clk, Q => 
                           n_1243, QN => n8854);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1720, CK => Clk, Q => 
                           n_1244, QN => n8855);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1719, CK => Clk, Q => 
                           n_1245, QN => n8856);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1718, CK => Clk, Q => 
                           n_1246, QN => n8857);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1789, CK => Clk, Q => 
                           n_1247, QN => n8786);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1788, CK => Clk, Q => 
                           n_1248, QN => n8787);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1787, CK => Clk, Q => 
                           n_1249, QN => n8788);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1786, CK => Clk, Q => 
                           n_1250, QN => n8789);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1785, CK => Clk, Q => 
                           n_1251, QN => n8790);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1784, CK => Clk, Q => 
                           n_1252, QN => n8791);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1783, CK => Clk, Q => 
                           n_1253, QN => n8792);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1782, CK => Clk, Q => 
                           n_1254, QN => n8793);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2173, CK => Clk, Q => 
                           n_1255, QN => n8402);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2172, CK => Clk, Q => 
                           n_1256, QN => n8403);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2171, CK => Clk, Q => 
                           n_1257, QN => n8404);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2170, CK => Clk, Q => 
                           n_1258, QN => n8405);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2169, CK => Clk, Q => 
                           n_1259, QN => n8406);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2168, CK => Clk, Q => 
                           n_1260, QN => n8407);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2167, CK => Clk, Q => 
                           n_1261, QN => n8408);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2166, CK => Clk, Q => 
                           n_1262, QN => n8409);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1917, CK => Clk, Q => 
                           n_1263, QN => n8658);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1916, CK => Clk, Q => 
                           n_1264, QN => n8659);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1915, CK => Clk, Q => 
                           n_1265, QN => n8660);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1914, CK => Clk, Q => 
                           n_1266, QN => n8661);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1913, CK => Clk, Q => 
                           n_1267, QN => n8662);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1912, CK => Clk, Q => 
                           n_1268, QN => n8663);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1911, CK => Clk, Q => 
                           n_1269, QN => n8664);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1910, CK => Clk, Q => 
                           n_1270, QN => n8665);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2141, CK => Clk, Q => 
                           n_1271, QN => n8434);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2140, CK => Clk, Q => 
                           n_1272, QN => n8435);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2139, CK => Clk, Q => 
                           n_1273, QN => n8436);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2138, CK => Clk, Q => 
                           n_1274, QN => n8437);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2137, CK => Clk, Q => 
                           n_1275, QN => n8438);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2136, CK => Clk, Q => 
                           n_1276, QN => n8439);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2135, CK => Clk, Q => 
                           n_1277, QN => n8440);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2134, CK => Clk, Q => 
                           n_1278, QN => n8441);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1333, CK => Clk, Q => 
                           n_1279, QN => n9242);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1332, CK => Clk, Q => 
                           n_1280, QN => n9243);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1331, CK => Clk, Q => 
                           n_1281, QN => n9244);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1330, CK => Clk, Q => 
                           n_1282, QN => n9245);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1329, CK => Clk, Q => 
                           n_1283, QN => n9246);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1328, CK => Clk, Q => 
                           n_1284, QN => n9247);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1327, CK => Clk, Q => 
                           n_1285, QN => n9248);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1326, CK => Clk, Q => 
                           n_1286, QN => n9249);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1325, CK => Clk, Q => 
                           n_1287, QN => n9250);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1324, CK => Clk, Q => 
                           n_1288, QN => n9251);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1323, CK => Clk, Q => 
                           n_1289, QN => n9252);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1322, CK => Clk, Q => 
                           n_1290, QN => n9253);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1321, CK => Clk, Q => 
                           n_1291, QN => n9254);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1320, CK => Clk, Q => 
                           n_1292, QN => n9255);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1319, CK => Clk, Q => 
                           n_1293, QN => n9256);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1318, CK => Clk, Q => 
                           n_1294, QN => n9257);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1317, CK => Clk, Q => 
                           n_1295, QN => n9258);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1316, CK => Clk, Q => 
                           n_1296, QN => n9259);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1315, CK => Clk, Q => 
                           n_1297, QN => n9260);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1314, CK => Clk, Q => 
                           n_1298, QN => n9261);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1313, CK => Clk, Q => 
                           n_1299, QN => n9262);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1312, CK => Clk, Q => 
                           n_1300, QN => n9263);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1311, CK => Clk, Q => 
                           n_1301, QN => n9264);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1310, CK => Clk, Q => 
                           n_1302, QN => n9265);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1493, CK => Clk, Q => 
                           n_1303, QN => n9082);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1492, CK => Clk, Q => 
                           n_1304, QN => n9083);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1491, CK => Clk, Q => 
                           n_1305, QN => n9084);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1490, CK => Clk, Q => 
                           n_1306, QN => n9085);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1489, CK => Clk, Q => 
                           n_1307, QN => n9086);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1488, CK => Clk, Q => 
                           n_1308, QN => n9087);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1487, CK => Clk, Q => 
                           n_1309, QN => n9088);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1486, CK => Clk, Q => 
                           n_1310, QN => n9089);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1485, CK => Clk, Q => 
                           n_1311, QN => n9090);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1484, CK => Clk, Q => 
                           n_1312, QN => n9091);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1483, CK => Clk, Q => 
                           n_1313, QN => n9092);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1482, CK => Clk, Q => 
                           n_1314, QN => n9093);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1481, CK => Clk, Q => 
                           n_1315, QN => n9094);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1480, CK => Clk, Q => 
                           n_1316, QN => n9095);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1479, CK => Clk, Q => 
                           n_1317, QN => n9096);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1478, CK => Clk, Q => 
                           n_1318, QN => n9097);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1477, CK => Clk, Q => 
                           n_1319, QN => n9098);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1476, CK => Clk, Q => 
                           n_1320, QN => n9099);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1475, CK => Clk, Q => 
                           n_1321, QN => n9100);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1474, CK => Clk, Q => 
                           n_1322, QN => n9101);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1473, CK => Clk, Q => 
                           n_1323, QN => n9102);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1472, CK => Clk, Q => 
                           n_1324, QN => n9103);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1471, CK => Clk, Q => 
                           n_1325, QN => n9104);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1470, CK => Clk, Q => 
                           n_1326, QN => n9105);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1621, CK => Clk, Q => 
                           n_1327, QN => n8954);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1620, CK => Clk, Q => 
                           n_1328, QN => n8955);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1619, CK => Clk, Q => 
                           n_1329, QN => n8956);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1618, CK => Clk, Q => 
                           n_1330, QN => n8957);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1617, CK => Clk, Q => 
                           n_1331, QN => n8958);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1616, CK => Clk, Q => 
                           n_1332, QN => n8959);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1615, CK => Clk, Q => 
                           n_1333, QN => n8960);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1614, CK => Clk, Q => 
                           n_1334, QN => n8961);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1613, CK => Clk, Q => 
                           n_1335, QN => n8962);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1612, CK => Clk, Q => 
                           n_1336, QN => n8963);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1611, CK => Clk, Q => 
                           n_1337, QN => n8964);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1610, CK => Clk, Q => 
                           n_1338, QN => n8965);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1609, CK => Clk, Q => 
                           n_1339, QN => n8966);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1608, CK => Clk, Q => 
                           n_1340, QN => n8967);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1607, CK => Clk, Q => 
                           n_1341, QN => n8968);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1606, CK => Clk, Q => 
                           n_1342, QN => n8969);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1605, CK => Clk, Q => 
                           n_1343, QN => n8970);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1604, CK => Clk, Q => 
                           n_1344, QN => n8971);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1603, CK => Clk, Q => 
                           n_1345, QN => n8972);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1602, CK => Clk, Q => 
                           n_1346, QN => n8973);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1601, CK => Clk, Q => 
                           n_1347, QN => n8974);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1600, CK => Clk, Q => 
                           n_1348, QN => n8975);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1599, CK => Clk, Q => 
                           n_1349, QN => n8976);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1598, CK => Clk, Q => 
                           n_1350, QN => n8977);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1653, CK => Clk, Q => 
                           n_1351, QN => n8922);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1652, CK => Clk, Q => 
                           n_1352, QN => n8923);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1651, CK => Clk, Q => 
                           n_1353, QN => n8924);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1650, CK => Clk, Q => 
                           n_1354, QN => n8925);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1649, CK => Clk, Q => 
                           n_1355, QN => n8926);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1648, CK => Clk, Q => 
                           n_1356, QN => n8927);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1647, CK => Clk, Q => 
                           n_1357, QN => n8928);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1646, CK => Clk, Q => 
                           n_1358, QN => n8929);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1645, CK => Clk, Q => 
                           n_1359, QN => n8930);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1644, CK => Clk, Q => 
                           n_1360, QN => n8931);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1643, CK => Clk, Q => 
                           n_1361, QN => n8932);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1642, CK => Clk, Q => 
                           n_1362, QN => n8933);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1641, CK => Clk, Q => 
                           n_1363, QN => n8934);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1640, CK => Clk, Q => 
                           n_1364, QN => n8935);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1639, CK => Clk, Q => 
                           n_1365, QN => n8936);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1638, CK => Clk, Q => 
                           n_1366, QN => n8937);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1637, CK => Clk, Q => 
                           n_1367, QN => n8938);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1636, CK => Clk, Q => 
                           n_1368, QN => n8939);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1635, CK => Clk, Q => 
                           n_1369, QN => n8940);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1634, CK => Clk, Q => 
                           n_1370, QN => n8941);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1633, CK => Clk, Q => 
                           n_1371, QN => n8942);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1632, CK => Clk, Q => 
                           n_1372, QN => n8943);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1631, CK => Clk, Q => 
                           n_1373, QN => n8944);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1630, CK => Clk, Q => 
                           n_1374, QN => n8945);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1941, CK => Clk, Q => 
                           n_1375, QN => n8634);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1940, CK => Clk, Q => 
                           n_1376, QN => n8635);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1939, CK => Clk, Q => 
                           n_1377, QN => n8636);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1938, CK => Clk, Q => 
                           n_1378, QN => n8637);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1937, CK => Clk, Q => 
                           n_1379, QN => n8638);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1936, CK => Clk, Q => 
                           n_1380, QN => n8639);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1935, CK => Clk, Q => 
                           n_1381, QN => n8640);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1934, CK => Clk, Q => 
                           n_1382, QN => n8641);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1933, CK => Clk, Q => 
                           n_1383, QN => n8642);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1932, CK => Clk, Q => 
                           n_1384, QN => n8643);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1931, CK => Clk, Q => 
                           n_1385, QN => n8644);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1930, CK => Clk, Q => 
                           n_1386, QN => n8645);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1929, CK => Clk, Q => 
                           n_1387, QN => n8646);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1928, CK => Clk, Q => 
                           n_1388, QN => n8647);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1927, CK => Clk, Q => 
                           n_1389, QN => n8648);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1926, CK => Clk, Q => 
                           n_1390, QN => n8649);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1925, CK => Clk, Q => 
                           n_1391, QN => n8650);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1924, CK => Clk, Q => 
                           n_1392, QN => n8651);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1923, CK => Clk, Q => 
                           n_1393, QN => n8652);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1922, CK => Clk, Q => 
                           n_1394, QN => n8653);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1921, CK => Clk, Q => 
                           n_1395, QN => n8654);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1920, CK => Clk, Q => 
                           n_1396, QN => n8655);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1919, CK => Clk, Q => 
                           n_1397, QN => n8656);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1918, CK => Clk, Q => 
                           n_1398, QN => n8657);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1877, CK => Clk, Q => 
                           n_1399, QN => n8698);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1876, CK => Clk, Q => 
                           n_1400, QN => n8699);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1875, CK => Clk, Q => 
                           n_1401, QN => n8700);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1874, CK => Clk, Q => 
                           n_1402, QN => n8701);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1873, CK => Clk, Q => 
                           n_1403, QN => n8702);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1872, CK => Clk, Q => 
                           n_1404, QN => n8703);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1871, CK => Clk, Q => 
                           n_1405, QN => n8704);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1870, CK => Clk, Q => 
                           n_1406, QN => n8705);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1869, CK => Clk, Q => 
                           n_1407, QN => n8706);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1868, CK => Clk, Q => 
                           n_1408, QN => n8707);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1867, CK => Clk, Q => 
                           n_1409, QN => n8708);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1866, CK => Clk, Q => 
                           n_1410, QN => n8709);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1865, CK => Clk, Q => 
                           n_1411, QN => n8710);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1864, CK => Clk, Q => 
                           n_1412, QN => n8711);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1863, CK => Clk, Q => 
                           n_1413, QN => n8712);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1862, CK => Clk, Q => 
                           n_1414, QN => n8713);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1861, CK => Clk, Q => 
                           n_1415, QN => n8714);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1860, CK => Clk, Q => 
                           n_1416, QN => n8715);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1859, CK => Clk, Q => 
                           n_1417, QN => n8716);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1858, CK => Clk, Q => 
                           n_1418, QN => n8717);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1857, CK => Clk, Q => 
                           n_1419, QN => n8718);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1856, CK => Clk, Q => 
                           n_1420, QN => n8719);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1855, CK => Clk, Q => 
                           n_1421, QN => n8720);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1854, CK => Clk, Q => 
                           n_1422, QN => n8721);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2229, CK => Clk, Q => 
                           n_1423, QN => n8346);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2228, CK => Clk, Q => 
                           n_1424, QN => n8347);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2227, CK => Clk, Q => 
                           n_1425, QN => n8348);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2226, CK => Clk, Q => 
                           n_1426, QN => n8349);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2225, CK => Clk, Q => 
                           n_1427, QN => n8350);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2224, CK => Clk, Q => 
                           n_1428, QN => n8351);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2223, CK => Clk, Q => 
                           n_1429, QN => n8352);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2222, CK => Clk, Q => 
                           n_1430, QN => n8353);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2221, CK => Clk, Q => 
                           n_1431, QN => n8354);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2220, CK => Clk, Q => 
                           n_1432, QN => n8355);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2219, CK => Clk, Q => 
                           n_1433, QN => n8356);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2218, CK => Clk, Q => 
                           n_1434, QN => n8357);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2217, CK => Clk, Q => 
                           n_1435, QN => n8358);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2216, CK => Clk, Q => 
                           n_1436, QN => n8359);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2215, CK => Clk, Q => n_1437
                           , QN => n8360);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2214, CK => Clk, Q => n_1438
                           , QN => n8361);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2213, CK => Clk, Q => n_1439
                           , QN => n8362);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2212, CK => Clk, Q => n_1440
                           , QN => n8363);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2211, CK => Clk, Q => n_1441
                           , QN => n8364);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2210, CK => Clk, Q => n_1442
                           , QN => n8365);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2209, CK => Clk, Q => n_1443
                           , QN => n8366);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2208, CK => Clk, Q => n_1444
                           , QN => n8367);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2207, CK => Clk, Q => n_1445
                           , QN => n8368);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2206, CK => Clk, Q => n_1446
                           , QN => n8369);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1365, CK => Clk, Q => 
                           n_1447, QN => n9210);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1364, CK => Clk, Q => 
                           n_1448, QN => n9211);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1363, CK => Clk, Q => 
                           n_1449, QN => n9212);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1362, CK => Clk, Q => 
                           n_1450, QN => n9213);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1361, CK => Clk, Q => 
                           n_1451, QN => n9214);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1360, CK => Clk, Q => 
                           n_1452, QN => n9215);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1359, CK => Clk, Q => 
                           n_1453, QN => n9216);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1358, CK => Clk, Q => 
                           n_1454, QN => n9217);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1357, CK => Clk, Q => 
                           n_1455, QN => n9218);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1356, CK => Clk, Q => 
                           n_1456, QN => n9219);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1355, CK => Clk, Q => 
                           n_1457, QN => n9220);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1354, CK => Clk, Q => 
                           n_1458, QN => n9221);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1353, CK => Clk, Q => 
                           n_1459, QN => n9222);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1352, CK => Clk, Q => 
                           n_1460, QN => n9223);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1351, CK => Clk, Q => 
                           n_1461, QN => n9224);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1350, CK => Clk, Q => 
                           n_1462, QN => n9225);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1349, CK => Clk, Q => 
                           n_1463, QN => n9226);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1348, CK => Clk, Q => 
                           n_1464, QN => n9227);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1347, CK => Clk, Q => 
                           n_1465, QN => n9228);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1346, CK => Clk, Q => 
                           n_1466, QN => n9229);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1345, CK => Clk, Q => 
                           n_1467, QN => n9230);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1344, CK => Clk, Q => 
                           n_1468, QN => n9231);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1343, CK => Clk, Q => 
                           n_1469, QN => n9232);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1342, CK => Clk, Q => 
                           n_1470, QN => n9233);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1397, CK => Clk, Q => 
                           n_1471, QN => n9178);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1396, CK => Clk, Q => 
                           n_1472, QN => n9179);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1395, CK => Clk, Q => 
                           n_1473, QN => n9180);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1394, CK => Clk, Q => 
                           n_1474, QN => n9181);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1393, CK => Clk, Q => 
                           n_1475, QN => n9182);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1392, CK => Clk, Q => 
                           n_1476, QN => n9183);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1391, CK => Clk, Q => 
                           n_1477, QN => n9184);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1390, CK => Clk, Q => 
                           n_1478, QN => n9185);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1389, CK => Clk, Q => 
                           n_1479, QN => n9186);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1388, CK => Clk, Q => 
                           n_1480, QN => n9187);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1387, CK => Clk, Q => 
                           n_1481, QN => n9188);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1386, CK => Clk, Q => 
                           n_1482, QN => n9189);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1385, CK => Clk, Q => 
                           n_1483, QN => n9190);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1384, CK => Clk, Q => 
                           n_1484, QN => n9191);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1383, CK => Clk, Q => 
                           n_1485, QN => n9192);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1382, CK => Clk, Q => 
                           n_1486, QN => n9193);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1381, CK => Clk, Q => 
                           n_1487, QN => n9194);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1380, CK => Clk, Q => 
                           n_1488, QN => n9195);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1379, CK => Clk, Q => 
                           n_1489, QN => n9196);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1378, CK => Clk, Q => 
                           n_1490, QN => n9197);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1377, CK => Clk, Q => 
                           n_1491, QN => n9198);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1376, CK => Clk, Q => 
                           n_1492, QN => n9199);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1375, CK => Clk, Q => 
                           n_1493, QN => n9200);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1374, CK => Clk, Q => 
                           n_1494, QN => n9201);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1685, CK => Clk, Q => 
                           n_1495, QN => n8890);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1684, CK => Clk, Q => 
                           n_1496, QN => n8891);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1683, CK => Clk, Q => 
                           n_1497, QN => n8892);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1682, CK => Clk, Q => 
                           n_1498, QN => n8893);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1681, CK => Clk, Q => 
                           n_1499, QN => n8894);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1680, CK => Clk, Q => 
                           n_1500, QN => n8895);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1679, CK => Clk, Q => 
                           n_1501, QN => n8896);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1678, CK => Clk, Q => 
                           n_1502, QN => n8897);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1677, CK => Clk, Q => 
                           n_1503, QN => n8898);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1676, CK => Clk, Q => 
                           n_1504, QN => n8899);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1675, CK => Clk, Q => 
                           n_1505, QN => n8900);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1674, CK => Clk, Q => 
                           n_1506, QN => n8901);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1673, CK => Clk, Q => 
                           n_1507, QN => n8902);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1672, CK => Clk, Q => 
                           n_1508, QN => n8903);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1671, CK => Clk, Q => 
                           n_1509, QN => n8904);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1670, CK => Clk, Q => 
                           n_1510, QN => n8905);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1669, CK => Clk, Q => 
                           n_1511, QN => n8906);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1668, CK => Clk, Q => 
                           n_1512, QN => n8907);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1667, CK => Clk, Q => 
                           n_1513, QN => n8908);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1666, CK => Clk, Q => 
                           n_1514, QN => n8909);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1665, CK => Clk, Q => 
                           n_1515, QN => n8910);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1664, CK => Clk, Q => 
                           n_1516, QN => n8911);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1663, CK => Clk, Q => 
                           n_1517, QN => n8912);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1662, CK => Clk, Q => 
                           n_1518, QN => n8913);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1717, CK => Clk, Q => 
                           n_1519, QN => n8858);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1716, CK => Clk, Q => 
                           n_1520, QN => n8859);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1715, CK => Clk, Q => 
                           n_1521, QN => n8860);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1714, CK => Clk, Q => 
                           n_1522, QN => n8861);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1713, CK => Clk, Q => 
                           n_1523, QN => n8862);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1712, CK => Clk, Q => 
                           n_1524, QN => n8863);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1711, CK => Clk, Q => 
                           n_1525, QN => n8864);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1710, CK => Clk, Q => 
                           n_1526, QN => n8865);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1709, CK => Clk, Q => 
                           n_1527, QN => n8866);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1708, CK => Clk, Q => 
                           n_1528, QN => n8867);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1707, CK => Clk, Q => 
                           n_1529, QN => n8868);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1706, CK => Clk, Q => 
                           n_1530, QN => n8869);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1705, CK => Clk, Q => 
                           n_1531, QN => n8870);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1704, CK => Clk, Q => 
                           n_1532, QN => n8871);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1703, CK => Clk, Q => 
                           n_1533, QN => n8872);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1702, CK => Clk, Q => 
                           n_1534, QN => n8873);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1701, CK => Clk, Q => 
                           n_1535, QN => n8874);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1700, CK => Clk, Q => 
                           n_1536, QN => n8875);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1699, CK => Clk, Q => 
                           n_1537, QN => n8876);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1698, CK => Clk, Q => 
                           n_1538, QN => n8877);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1697, CK => Clk, Q => 
                           n_1539, QN => n8878);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1696, CK => Clk, Q => 
                           n_1540, QN => n8879);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1695, CK => Clk, Q => 
                           n_1541, QN => n8880);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1694, CK => Clk, Q => 
                           n_1542, QN => n8881);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1781, CK => Clk, Q => 
                           n_1543, QN => n8794);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1780, CK => Clk, Q => 
                           n_1544, QN => n8795);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1779, CK => Clk, Q => 
                           n_1545, QN => n8796);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1778, CK => Clk, Q => 
                           n_1546, QN => n8797);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1777, CK => Clk, Q => 
                           n_1547, QN => n8798);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1776, CK => Clk, Q => 
                           n_1548, QN => n8799);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1775, CK => Clk, Q => 
                           n_1549, QN => n8800);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1774, CK => Clk, Q => 
                           n_1550, QN => n8801);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1773, CK => Clk, Q => 
                           n_1551, QN => n8802);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1772, CK => Clk, Q => 
                           n_1552, QN => n8803);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1771, CK => Clk, Q => 
                           n_1553, QN => n8804);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1770, CK => Clk, Q => 
                           n_1554, QN => n8805);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1769, CK => Clk, Q => 
                           n_1555, QN => n8806);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1768, CK => Clk, Q => 
                           n_1556, QN => n8807);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1767, CK => Clk, Q => 
                           n_1557, QN => n8808);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1766, CK => Clk, Q => 
                           n_1558, QN => n8809);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1765, CK => Clk, Q => 
                           n_1559, QN => n8810);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1764, CK => Clk, Q => 
                           n_1560, QN => n8811);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1763, CK => Clk, Q => 
                           n_1561, QN => n8812);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1762, CK => Clk, Q => 
                           n_1562, QN => n8813);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1761, CK => Clk, Q => 
                           n_1563, QN => n8814);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1760, CK => Clk, Q => 
                           n_1564, QN => n8815);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1759, CK => Clk, Q => 
                           n_1565, QN => n8816);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1758, CK => Clk, Q => 
                           n_1566, QN => n8817);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2165, CK => Clk, Q => 
                           n_1567, QN => n8410);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2164, CK => Clk, Q => 
                           n_1568, QN => n8411);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2163, CK => Clk, Q => 
                           n_1569, QN => n8412);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2162, CK => Clk, Q => 
                           n_1570, QN => n8413);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2161, CK => Clk, Q => 
                           n_1571, QN => n8414);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2160, CK => Clk, Q => 
                           n_1572, QN => n8415);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2159, CK => Clk, Q => 
                           n_1573, QN => n8416);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2158, CK => Clk, Q => 
                           n_1574, QN => n8417);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2157, CK => Clk, Q => 
                           n_1575, QN => n8418);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2156, CK => Clk, Q => 
                           n_1576, QN => n8419);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2155, CK => Clk, Q => 
                           n_1577, QN => n8420);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2154, CK => Clk, Q => 
                           n_1578, QN => n8421);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2153, CK => Clk, Q => 
                           n_1579, QN => n8422);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2152, CK => Clk, Q => 
                           n_1580, QN => n8423);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2151, CK => Clk, Q => n_1581
                           , QN => n8424);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2150, CK => Clk, Q => n_1582
                           , QN => n8425);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2149, CK => Clk, Q => n_1583
                           , QN => n8426);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2148, CK => Clk, Q => n_1584
                           , QN => n8427);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2147, CK => Clk, Q => n_1585
                           , QN => n8428);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2146, CK => Clk, Q => n_1586
                           , QN => n8429);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2145, CK => Clk, Q => n_1587
                           , QN => n8430);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2144, CK => Clk, Q => n_1588
                           , QN => n8431);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2143, CK => Clk, Q => n_1589
                           , QN => n8432);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2142, CK => Clk, Q => n_1590
                           , QN => n8433);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1909, CK => Clk, Q => 
                           n_1591, QN => n8666);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1908, CK => Clk, Q => 
                           n_1592, QN => n8667);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1907, CK => Clk, Q => 
                           n_1593, QN => n8668);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1906, CK => Clk, Q => 
                           n_1594, QN => n8669);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1905, CK => Clk, Q => 
                           n_1595, QN => n8670);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1904, CK => Clk, Q => 
                           n_1596, QN => n8671);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1903, CK => Clk, Q => 
                           n_1597, QN => n8672);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1902, CK => Clk, Q => 
                           n_1598, QN => n8673);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1901, CK => Clk, Q => 
                           n_1599, QN => n8674);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1900, CK => Clk, Q => 
                           n_1600, QN => n8675);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1899, CK => Clk, Q => 
                           n_1601, QN => n8676);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1898, CK => Clk, Q => 
                           n_1602, QN => n8677);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1897, CK => Clk, Q => 
                           n_1603, QN => n8678);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1896, CK => Clk, Q => 
                           n_1604, QN => n8679);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1895, CK => Clk, Q => 
                           n_1605, QN => n8680);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1894, CK => Clk, Q => 
                           n_1606, QN => n8681);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1893, CK => Clk, Q => 
                           n_1607, QN => n8682);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1892, CK => Clk, Q => 
                           n_1608, QN => n8683);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1891, CK => Clk, Q => 
                           n_1609, QN => n8684);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1890, CK => Clk, Q => 
                           n_1610, QN => n8685);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1889, CK => Clk, Q => 
                           n_1611, QN => n8686);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1888, CK => Clk, Q => 
                           n_1612, QN => n8687);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1887, CK => Clk, Q => 
                           n_1613, QN => n8688);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1886, CK => Clk, Q => 
                           n_1614, QN => n8689);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2133, CK => Clk, Q => 
                           n_1615, QN => n8442);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2132, CK => Clk, Q => 
                           n_1616, QN => n8443);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2131, CK => Clk, Q => 
                           n_1617, QN => n8444);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2130, CK => Clk, Q => 
                           n_1618, QN => n8445);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2129, CK => Clk, Q => 
                           n_1619, QN => n8446);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2128, CK => Clk, Q => 
                           n_1620, QN => n8447);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2127, CK => Clk, Q => 
                           n_1621, QN => n8448);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2126, CK => Clk, Q => 
                           n_1622, QN => n8449);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2125, CK => Clk, Q => 
                           n_1623, QN => n8450);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2124, CK => Clk, Q => 
                           n_1624, QN => n8451);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2123, CK => Clk, Q => 
                           n_1625, QN => n8452);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2122, CK => Clk, Q => 
                           n_1626, QN => n8453);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2121, CK => Clk, Q => 
                           n_1627, QN => n8454);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2120, CK => Clk, Q => 
                           n_1628, QN => n8455);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2119, CK => Clk, Q => n_1629
                           , QN => n8456);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2118, CK => Clk, Q => n_1630
                           , QN => n8457);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2117, CK => Clk, Q => n_1631
                           , QN => n8458);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2116, CK => Clk, Q => n_1632
                           , QN => n8459);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2115, CK => Clk, Q => n_1633
                           , QN => n8460);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2114, CK => Clk, Q => n_1634
                           , QN => n8461);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2113, CK => Clk, Q => n_1635
                           , QN => n8462);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2112, CK => Clk, Q => n_1636
                           , QN => n8463);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2111, CK => Clk, Q => n_1637
                           , QN => n8464);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2110, CK => Clk, Q => n_1638
                           , QN => n8465);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1469, CK => Clk, Q => 
                           n7396, QN => n9106);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1468, CK => Clk, Q => 
                           n7395, QN => n9107);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1467, CK => Clk, Q => 
                           n7394, QN => n9108);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1466, CK => Clk, Q => 
                           n7393, QN => n9109);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1465, CK => Clk, Q => 
                           n7392, QN => n9110);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1464, CK => Clk, Q => 
                           n7391, QN => n9111);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1463, CK => Clk, Q => 
                           n7390, QN => n9112);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1462, CK => Clk, Q => 
                           n7389, QN => n9113);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1597, CK => Clk, Q => 
                           n7588, QN => n8978);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1596, CK => Clk, Q => 
                           n7587, QN => n8979);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1595, CK => Clk, Q => 
                           n7586, QN => n8980);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1594, CK => Clk, Q => 
                           n7585, QN => n8981);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1593, CK => Clk, Q => 
                           n7584, QN => n8982);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1592, CK => Clk, Q => 
                           n7583, QN => n8983);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1591, CK => Clk, Q => 
                           n7582, QN => n8984);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1590, CK => Clk, Q => 
                           n7581, QN => n8985);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1757, CK => Clk, Q => 
                           n7492, QN => n8818);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1756, CK => Clk, Q => 
                           n7491, QN => n8819);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1755, CK => Clk, Q => 
                           n7490, QN => n8820);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1754, CK => Clk, Q => 
                           n7489, QN => n8821);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1753, CK => Clk, Q => 
                           n7488, QN => n8822);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1752, CK => Clk, Q => 
                           n7487, QN => n8823);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1751, CK => Clk, Q => 
                           n7486, QN => n8824);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1750, CK => Clk, Q => 
                           n7485, QN => n8825);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1821, CK => Clk, Q => 
                           n11004, QN => n8754);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1820, CK => Clk, Q => 
                           n11003, QN => n8755);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1819, CK => Clk, Q => 
                           n11002, QN => n8756);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1818, CK => Clk, Q => 
                           n11001, QN => n8757);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1817, CK => Clk, Q => 
                           n11000, QN => n8758);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1816, CK => Clk, Q => 
                           n10999, QN => n8759);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1815, CK => Clk, Q => 
                           n10998, QN => n8760);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1814, CK => Clk, Q => 
                           n10997, QN => n8761);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2013, CK => Clk, Q => 
                           n10716, QN => n8562);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2012, CK => Clk, Q => 
                           n10715, QN => n8563);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2011, CK => Clk, Q => 
                           n10714, QN => n8564);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2010, CK => Clk, Q => 
                           n10713, QN => n8565);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2009, CK => Clk, Q => 
                           n10712, QN => n8566);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2008, CK => Clk, Q => 
                           n10711, QN => n8567);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2007, CK => Clk, Q => 
                           n10710, QN => n8568);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2006, CK => Clk, Q => 
                           n10709, QN => n8569);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2109, CK => Clk, Q => 
                           n11164, QN => n8466);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2108, CK => Clk, Q => 
                           n11163, QN => n8467);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2107, CK => Clk, Q => 
                           n11162, QN => n8468);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2106, CK => Clk, Q => 
                           n11161, QN => n8469);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2105, CK => Clk, Q => 
                           n11160, QN => n8470);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2104, CK => Clk, Q => 
                           n11159, QN => n8471);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2103, CK => Clk, Q => 
                           n11158, QN => n8472);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2102, CK => Clk, Q => 
                           n11157, QN => n8473);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2301, CK => Clk, Q => 
                           n10876, QN => n8274);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2300, CK => Clk, Q => 
                           n10875, QN => n8275);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2299, CK => Clk, Q => 
                           n10874, QN => n8276);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2298, CK => Clk, Q => 
                           n10873, QN => n8277);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2297, CK => Clk, Q => 
                           n10872, QN => n8278);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2296, CK => Clk, Q => 
                           n10871, QN => n8279);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2295, CK => Clk, Q => 
                           n10870, QN => n8280);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2294, CK => Clk, Q => 
                           n10869, QN => n8281);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1461, CK => Clk, Q => 
                           n7388, QN => n9114);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1460, CK => Clk, Q => 
                           n7387, QN => n9115);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1459, CK => Clk, Q => 
                           n7386, QN => n9116);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1458, CK => Clk, Q => 
                           n7385, QN => n9117);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1457, CK => Clk, Q => 
                           n7384, QN => n9118);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1456, CK => Clk, Q => 
                           n7383, QN => n9119);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1455, CK => Clk, Q => 
                           n7382, QN => n9120);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1454, CK => Clk, Q => 
                           n7381, QN => n9121);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1453, CK => Clk, Q => 
                           n7380, QN => n9122);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1452, CK => Clk, Q => 
                           n7379, QN => n9123);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1451, CK => Clk, Q => 
                           n7378, QN => n9124);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1450, CK => Clk, Q => 
                           n7377, QN => n9125);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1449, CK => Clk, Q => 
                           n7376, QN => n9126);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1448, CK => Clk, Q => 
                           n7375, QN => n9127);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1447, CK => Clk, Q => n7374
                           , QN => n9128);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1446, CK => Clk, Q => n7397
                           , QN => n9129);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1445, CK => Clk, Q => n7405
                           , QN => n9130);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1444, CK => Clk, Q => n7404
                           , QN => n9131);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1443, CK => Clk, Q => n7403
                           , QN => n9132);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1442, CK => Clk, Q => n7402
                           , QN => n9133);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1441, CK => Clk, Q => n7401
                           , QN => n9134);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1440, CK => Clk, Q => n7400
                           , QN => n9135);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1439, CK => Clk, Q => n7399
                           , QN => n9136);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1438, CK => Clk, Q => n7398
                           , QN => n9137);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1589, CK => Clk, Q => 
                           n7580, QN => n8986);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1588, CK => Clk, Q => 
                           n7579, QN => n8987);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1587, CK => Clk, Q => 
                           n7578, QN => n8988);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1586, CK => Clk, Q => 
                           n7577, QN => n8989);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1585, CK => Clk, Q => 
                           n7576, QN => n8990);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1584, CK => Clk, Q => 
                           n7575, QN => n8991);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1583, CK => Clk, Q => 
                           n7574, QN => n8992);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1582, CK => Clk, Q => 
                           n7573, QN => n8993);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1581, CK => Clk, Q => 
                           n7572, QN => n8994);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1580, CK => Clk, Q => 
                           n7571, QN => n8995);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1579, CK => Clk, Q => 
                           n7570, QN => n8996);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1578, CK => Clk, Q => 
                           n7569, QN => n8997);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1577, CK => Clk, Q => 
                           n7568, QN => n8998);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1576, CK => Clk, Q => 
                           n7567, QN => n8999);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1575, CK => Clk, Q => n7566
                           , QN => n9000);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1574, CK => Clk, Q => n7589
                           , QN => n9001);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1573, CK => Clk, Q => n7597
                           , QN => n9002);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1572, CK => Clk, Q => n7596
                           , QN => n9003);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1571, CK => Clk, Q => n7595
                           , QN => n9004);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1570, CK => Clk, Q => n7594
                           , QN => n9005);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1569, CK => Clk, Q => n7593
                           , QN => n9006);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1568, CK => Clk, Q => n7592
                           , QN => n9007);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1567, CK => Clk, Q => n7591
                           , QN => n9008);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1566, CK => Clk, Q => n7590
                           , QN => n9009);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1749, CK => Clk, Q => 
                           n7484, QN => n8826);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1748, CK => Clk, Q => 
                           n7483, QN => n8827);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1747, CK => Clk, Q => 
                           n7482, QN => n8828);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1746, CK => Clk, Q => 
                           n7481, QN => n8829);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1745, CK => Clk, Q => 
                           n7480, QN => n8830);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1744, CK => Clk, Q => 
                           n7479, QN => n8831);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1743, CK => Clk, Q => 
                           n7478, QN => n8832);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1742, CK => Clk, Q => 
                           n7477, QN => n8833);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1741, CK => Clk, Q => 
                           n7476, QN => n8834);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1740, CK => Clk, Q => 
                           n7475, QN => n8835);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1739, CK => Clk, Q => 
                           n7474, QN => n8836);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1738, CK => Clk, Q => 
                           n7473, QN => n8837);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1737, CK => Clk, Q => 
                           n7472, QN => n8838);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1736, CK => Clk, Q => 
                           n7471, QN => n8839);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1735, CK => Clk, Q => n7470
                           , QN => n8840);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1734, CK => Clk, Q => n7493
                           , QN => n8841);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1733, CK => Clk, Q => n7501
                           , QN => n8842);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1732, CK => Clk, Q => n7500
                           , QN => n8843);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1731, CK => Clk, Q => n7499
                           , QN => n8844);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1730, CK => Clk, Q => n7498
                           , QN => n8845);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1729, CK => Clk, Q => n7497
                           , QN => n8846);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1728, CK => Clk, Q => n7496
                           , QN => n8847);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1727, CK => Clk, Q => n7495
                           , QN => n8848);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1726, CK => Clk, Q => n7494
                           , QN => n8849);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1813, CK => Clk, Q => 
                           n10996, QN => n8762);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1812, CK => Clk, Q => 
                           n10995, QN => n8763);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1811, CK => Clk, Q => 
                           n10994, QN => n8764);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1810, CK => Clk, Q => 
                           n10993, QN => n8765);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1809, CK => Clk, Q => 
                           n10992, QN => n8766);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1808, CK => Clk, Q => 
                           n10991, QN => n8767);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1807, CK => Clk, Q => 
                           n10990, QN => n8768);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1806, CK => Clk, Q => 
                           n10989, QN => n8769);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1805, CK => Clk, Q => 
                           n10988, QN => n8770);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1804, CK => Clk, Q => 
                           n10987, QN => n8771);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1803, CK => Clk, Q => 
                           n10986, QN => n8772);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1802, CK => Clk, Q => 
                           n10985, QN => n8773);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1801, CK => Clk, Q => 
                           n10984, QN => n8774);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1800, CK => Clk, Q => 
                           n10983, QN => n8775);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1799, CK => Clk, Q => 
                           n10982, QN => n8776);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1798, CK => Clk, Q => 
                           n10981, QN => n8777);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1797, CK => Clk, Q => 
                           n10980, QN => n8778);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1796, CK => Clk, Q => 
                           n10979, QN => n8779);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1795, CK => Clk, Q => 
                           n10978, QN => n8780);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1794, CK => Clk, Q => 
                           n10977, QN => n8781);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1793, CK => Clk, Q => 
                           n10976, QN => n8782);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1792, CK => Clk, Q => 
                           n10975, QN => n8783);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1791, CK => Clk, Q => 
                           n10974, QN => n8784);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1790, CK => Clk, Q => 
                           n10973, QN => n8785);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2005, CK => Clk, Q => 
                           n10708, QN => n8570);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2004, CK => Clk, Q => 
                           n10707, QN => n8571);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2003, CK => Clk, Q => 
                           n10706, QN => n8572);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2002, CK => Clk, Q => 
                           n10705, QN => n8573);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2001, CK => Clk, Q => 
                           n10704, QN => n8574);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2000, CK => Clk, Q => 
                           n10703, QN => n8575);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1999, CK => Clk, Q => 
                           n10702, QN => n8576);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1998, CK => Clk, Q => 
                           n10701, QN => n8577);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1997, CK => Clk, Q => 
                           n10700, QN => n8578);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1996, CK => Clk, Q => 
                           n10699, QN => n8579);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1995, CK => Clk, Q => 
                           n10698, QN => n8580);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1994, CK => Clk, Q => 
                           n10697, QN => n8581);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1993, CK => Clk, Q => 
                           n10696, QN => n8582);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1992, CK => Clk, Q => 
                           n10695, QN => n8583);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1991, CK => Clk, Q => n10694
                           , QN => n8584);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1990, CK => Clk, Q => n10693
                           , QN => n8585);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1989, CK => Clk, Q => n10692
                           , QN => n8586);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1988, CK => Clk, Q => n10691
                           , QN => n8587);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1987, CK => Clk, Q => n10690
                           , QN => n8588);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1986, CK => Clk, Q => n10689
                           , QN => n8589);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1985, CK => Clk, Q => n10688
                           , QN => n8590);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1984, CK => Clk, Q => n10687
                           , QN => n8591);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1983, CK => Clk, Q => n10686
                           , QN => n8592);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1982, CK => Clk, Q => n10685
                           , QN => n8593);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2101, CK => Clk, Q => 
                           n11156, QN => n8474);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2100, CK => Clk, Q => 
                           n11155, QN => n8475);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2099, CK => Clk, Q => 
                           n11154, QN => n8476);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2098, CK => Clk, Q => 
                           n11153, QN => n8477);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2097, CK => Clk, Q => 
                           n11152, QN => n8478);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2096, CK => Clk, Q => 
                           n11151, QN => n8479);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2095, CK => Clk, Q => 
                           n11150, QN => n8480);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2094, CK => Clk, Q => 
                           n11149, QN => n8481);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2093, CK => Clk, Q => 
                           n11148, QN => n8482);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2092, CK => Clk, Q => 
                           n11147, QN => n8483);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2091, CK => Clk, Q => 
                           n11146, QN => n8484);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2090, CK => Clk, Q => 
                           n11145, QN => n8485);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2089, CK => Clk, Q => 
                           n11144, QN => n8486);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2088, CK => Clk, Q => 
                           n11143, QN => n8487);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2087, CK => Clk, Q => n11142
                           , QN => n8488);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2086, CK => Clk, Q => n11141
                           , QN => n8489);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2085, CK => Clk, Q => n11140
                           , QN => n8490);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2084, CK => Clk, Q => n11139
                           , QN => n8491);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2083, CK => Clk, Q => n11138
                           , QN => n8492);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2082, CK => Clk, Q => n11137
                           , QN => n8493);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2081, CK => Clk, Q => n11136
                           , QN => n8494);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2080, CK => Clk, Q => n11135
                           , QN => n8495);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2079, CK => Clk, Q => n11134
                           , QN => n8496);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2078, CK => Clk, Q => n11133
                           , QN => n8497);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2293, CK => Clk, Q => 
                           n10868, QN => n8282);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2292, CK => Clk, Q => 
                           n10867, QN => n8283);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2291, CK => Clk, Q => 
                           n10866, QN => n8284);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2290, CK => Clk, Q => 
                           n10865, QN => n8285);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2289, CK => Clk, Q => 
                           n10864, QN => n8286);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2288, CK => Clk, Q => 
                           n10863, QN => n8287);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2287, CK => Clk, Q => 
                           n10862, QN => n8288);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2286, CK => Clk, Q => 
                           n10861, QN => n8289);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2285, CK => Clk, Q => 
                           n10860, QN => n8290);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2284, CK => Clk, Q => 
                           n10859, QN => n8291);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2283, CK => Clk, Q => 
                           n10858, QN => n8292);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2282, CK => Clk, Q => 
                           n10857, QN => n8293);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2281, CK => Clk, Q => 
                           n10856, QN => n8294);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2280, CK => Clk, Q => 
                           n10855, QN => n8295);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2279, CK => Clk, Q => n10854
                           , QN => n8296);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2278, CK => Clk, Q => n10853
                           , QN => n8297);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2277, CK => Clk, Q => n10852
                           , QN => n8298);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2276, CK => Clk, Q => n10851
                           , QN => n8299);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2275, CK => Clk, Q => n10850
                           , QN => n8300);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2274, CK => Clk, Q => n10849
                           , QN => n8301);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2273, CK => Clk, Q => n10848
                           , QN => n8302);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2272, CK => Clk, Q => n10847
                           , QN => n8303);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2271, CK => Clk, Q => n10846
                           , QN => n8304);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2270, CK => Clk, Q => n10845
                           , QN => n8305);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1437, CK => Clk, Q => 
                           n10940, QN => n9138);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1436, CK => Clk, Q => 
                           n10939, QN => n9139);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1435, CK => Clk, Q => 
                           n10938, QN => n9140);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1434, CK => Clk, Q => 
                           n10937, QN => n9141);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1433, CK => Clk, Q => 
                           n10936, QN => n9142);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1432, CK => Clk, Q => 
                           n10935, QN => n9143);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1431, CK => Clk, Q => 
                           n10934, QN => n9144);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1430, CK => Clk, Q => 
                           n10933, QN => n9145);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1533, CK => Clk, Q => 
                           n7556, QN => n9042);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1532, CK => Clk, Q => 
                           n7555, QN => n9043);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1531, CK => Clk, Q => 
                           n7554, QN => n9044);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1530, CK => Clk, Q => 
                           n7553, QN => n9045);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1529, CK => Clk, Q => 
                           n7552, QN => n9046);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1528, CK => Clk, Q => 
                           n7551, QN => n9047);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1527, CK => Clk, Q => 
                           n7550, QN => n9048);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1526, CK => Clk, Q => 
                           n7549, QN => n9049);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1565, CK => Clk, Q => 
                           n10972, QN => n9010);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1564, CK => Clk, Q => 
                           n10971, QN => n9011);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1563, CK => Clk, Q => 
                           n10970, QN => n9012);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1562, CK => Clk, Q => 
                           n10969, QN => n9013);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1561, CK => Clk, Q => 
                           n10968, QN => n9014);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1560, CK => Clk, Q => 
                           n10967, QN => n9015);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1559, CK => Clk, Q => 
                           n10966, QN => n9016);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1558, CK => Clk, Q => 
                           n10965, QN => n9017);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1853, CK => Clk, Q => 
                           n11036, QN => n8722);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1852, CK => Clk, Q => 
                           n11035, QN => n8723);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1851, CK => Clk, Q => 
                           n11034, QN => n8724);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1850, CK => Clk, Q => 
                           n11033, QN => n8725);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1849, CK => Clk, Q => 
                           n11032, QN => n8726);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1848, CK => Clk, Q => 
                           n11031, QN => n8727);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1847, CK => Clk, Q => 
                           n11030, QN => n8728);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1846, CK => Clk, Q => 
                           n11029, QN => n8729);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2045, CK => Clk, Q => 
                           n10748, QN => n8530);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2044, CK => Clk, Q => 
                           n10747, QN => n8531);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2043, CK => Clk, Q => 
                           n10746, QN => n8532);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2042, CK => Clk, Q => 
                           n10745, QN => n8533);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2041, CK => Clk, Q => 
                           n10744, QN => n8534);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2040, CK => Clk, Q => 
                           n10743, QN => n8535);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2039, CK => Clk, Q => 
                           n10742, QN => n8536);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2038, CK => Clk, Q => 
                           n10741, QN => n8537);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2077, CK => Clk, Q => 
                           n11132, QN => n8498);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2076, CK => Clk, Q => 
                           n11131, QN => n8499);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2075, CK => Clk, Q => 
                           n11130, QN => n8500);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2074, CK => Clk, Q => 
                           n11129, QN => n8501);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2073, CK => Clk, Q => 
                           n11128, QN => n8502);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2072, CK => Clk, Q => 
                           n11127, QN => n8503);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2071, CK => Clk, Q => 
                           n11126, QN => n8504);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2070, CK => Clk, Q => 
                           n11125, QN => n8505);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2205, CK => Clk, Q => 
                           n11196, QN => n8370);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2204, CK => Clk, Q => 
                           n11195, QN => n8371);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2203, CK => Clk, Q => 
                           n11194, QN => n8372);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2202, CK => Clk, Q => 
                           n11193, QN => n8373);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2201, CK => Clk, Q => 
                           n11192, QN => n8374);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2200, CK => Clk, Q => 
                           n11191, QN => n8375);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2199, CK => Clk, Q => 
                           n11190, QN => n8376);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2198, CK => Clk, Q => 
                           n11189, QN => n8377);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1429, CK => Clk, Q => 
                           n10932, QN => n9146);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1428, CK => Clk, Q => 
                           n10931, QN => n9147);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1427, CK => Clk, Q => 
                           n10930, QN => n9148);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1426, CK => Clk, Q => 
                           n10929, QN => n9149);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1425, CK => Clk, Q => 
                           n10928, QN => n9150);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1424, CK => Clk, Q => 
                           n10927, QN => n9151);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1423, CK => Clk, Q => 
                           n10926, QN => n9152);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1422, CK => Clk, Q => 
                           n10925, QN => n9153);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1421, CK => Clk, Q => 
                           n10924, QN => n9154);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1420, CK => Clk, Q => 
                           n10923, QN => n9155);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1419, CK => Clk, Q => 
                           n10922, QN => n9156);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1418, CK => Clk, Q => 
                           n10921, QN => n9157);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1417, CK => Clk, Q => 
                           n10920, QN => n9158);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1416, CK => Clk, Q => 
                           n10919, QN => n9159);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1415, CK => Clk, Q => 
                           n10918, QN => n9160);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1414, CK => Clk, Q => 
                           n10917, QN => n9161);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1413, CK => Clk, Q => 
                           n10916, QN => n9162);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1412, CK => Clk, Q => 
                           n10915, QN => n9163);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1411, CK => Clk, Q => 
                           n10914, QN => n9164);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1410, CK => Clk, Q => 
                           n10913, QN => n9165);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1409, CK => Clk, Q => 
                           n10912, QN => n9166);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1408, CK => Clk, Q => 
                           n10911, QN => n9167);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1407, CK => Clk, Q => 
                           n10910, QN => n9168);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1406, CK => Clk, Q => 
                           n10909, QN => n9169);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1525, CK => Clk, Q => 
                           n7548, QN => n9050);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1524, CK => Clk, Q => 
                           n7547, QN => n9051);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1523, CK => Clk, Q => 
                           n7546, QN => n9052);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1522, CK => Clk, Q => 
                           n7545, QN => n9053);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1521, CK => Clk, Q => 
                           n7544, QN => n9054);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1520, CK => Clk, Q => 
                           n7543, QN => n9055);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1519, CK => Clk, Q => 
                           n7542, QN => n9056);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1518, CK => Clk, Q => 
                           n7541, QN => n9057);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1517, CK => Clk, Q => 
                           n7540, QN => n9058);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1516, CK => Clk, Q => 
                           n7539, QN => n9059);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1515, CK => Clk, Q => 
                           n7538, QN => n9060);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1514, CK => Clk, Q => 
                           n7537, QN => n9061);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1513, CK => Clk, Q => 
                           n7536, QN => n9062);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1512, CK => Clk, Q => 
                           n7535, QN => n9063);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1511, CK => Clk, Q => n7534
                           , QN => n9064);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1510, CK => Clk, Q => n7557
                           , QN => n9065);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1509, CK => Clk, Q => n7565
                           , QN => n9066);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1508, CK => Clk, Q => n7564
                           , QN => n9067);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1507, CK => Clk, Q => n7563
                           , QN => n9068);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1506, CK => Clk, Q => n7562
                           , QN => n9069);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1505, CK => Clk, Q => n7561
                           , QN => n9070);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1504, CK => Clk, Q => n7560
                           , QN => n9071);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1503, CK => Clk, Q => n7559
                           , QN => n9072);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1502, CK => Clk, Q => n7558
                           , QN => n9073);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1557, CK => Clk, Q => 
                           n10964, QN => n9018);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1556, CK => Clk, Q => 
                           n10963, QN => n9019);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1555, CK => Clk, Q => 
                           n10962, QN => n9020);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1554, CK => Clk, Q => 
                           n10961, QN => n9021);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1553, CK => Clk, Q => 
                           n10960, QN => n9022);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1552, CK => Clk, Q => 
                           n10959, QN => n9023);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1551, CK => Clk, Q => 
                           n10958, QN => n9024);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1550, CK => Clk, Q => 
                           n10957, QN => n9025);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1549, CK => Clk, Q => 
                           n10956, QN => n9026);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1548, CK => Clk, Q => 
                           n10955, QN => n9027);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1547, CK => Clk, Q => 
                           n10954, QN => n9028);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1546, CK => Clk, Q => 
                           n10953, QN => n9029);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1545, CK => Clk, Q => 
                           n10952, QN => n9030);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1544, CK => Clk, Q => 
                           n10951, QN => n9031);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1543, CK => Clk, Q => 
                           n10950, QN => n9032);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1542, CK => Clk, Q => 
                           n10949, QN => n9033);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1541, CK => Clk, Q => 
                           n10948, QN => n9034);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1540, CK => Clk, Q => 
                           n10947, QN => n9035);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1539, CK => Clk, Q => 
                           n10946, QN => n9036);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1538, CK => Clk, Q => 
                           n10945, QN => n9037);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1537, CK => Clk, Q => 
                           n10944, QN => n9038);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1536, CK => Clk, Q => 
                           n10943, QN => n9039);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1535, CK => Clk, Q => 
                           n10942, QN => n9040);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1534, CK => Clk, Q => 
                           n10941, QN => n9041);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1845, CK => Clk, Q => 
                           n11028, QN => n8730);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1844, CK => Clk, Q => 
                           n11027, QN => n8731);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1843, CK => Clk, Q => 
                           n11026, QN => n8732);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1842, CK => Clk, Q => 
                           n11025, QN => n8733);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1841, CK => Clk, Q => 
                           n11024, QN => n8734);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1840, CK => Clk, Q => 
                           n11023, QN => n8735);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1839, CK => Clk, Q => 
                           n11022, QN => n8736);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1838, CK => Clk, Q => 
                           n11021, QN => n8737);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1837, CK => Clk, Q => 
                           n11020, QN => n8738);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1836, CK => Clk, Q => 
                           n11019, QN => n8739);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1835, CK => Clk, Q => 
                           n11018, QN => n8740);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1834, CK => Clk, Q => 
                           n11017, QN => n8741);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1833, CK => Clk, Q => 
                           n11016, QN => n8742);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1832, CK => Clk, Q => 
                           n11015, QN => n8743);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1831, CK => Clk, Q => 
                           n11014, QN => n8744);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1830, CK => Clk, Q => 
                           n11013, QN => n8745);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1829, CK => Clk, Q => 
                           n11012, QN => n8746);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1828, CK => Clk, Q => 
                           n11011, QN => n8747);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1827, CK => Clk, Q => 
                           n11010, QN => n8748);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1826, CK => Clk, Q => 
                           n11009, QN => n8749);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1825, CK => Clk, Q => 
                           n11008, QN => n8750);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1824, CK => Clk, Q => 
                           n11007, QN => n8751);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1823, CK => Clk, Q => 
                           n11006, QN => n8752);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1822, CK => Clk, Q => 
                           n11005, QN => n8753);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2037, CK => Clk, Q => 
                           n10740, QN => n8538);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2036, CK => Clk, Q => 
                           n10739, QN => n8539);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2035, CK => Clk, Q => 
                           n10738, QN => n8540);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2034, CK => Clk, Q => 
                           n10737, QN => n8541);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2033, CK => Clk, Q => 
                           n10736, QN => n8542);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2032, CK => Clk, Q => 
                           n10735, QN => n8543);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2031, CK => Clk, Q => 
                           n10734, QN => n8544);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2030, CK => Clk, Q => 
                           n10733, QN => n8545);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2029, CK => Clk, Q => 
                           n10732, QN => n8546);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2028, CK => Clk, Q => 
                           n10731, QN => n8547);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2027, CK => Clk, Q => 
                           n10730, QN => n8548);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2026, CK => Clk, Q => 
                           n10729, QN => n8549);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2025, CK => Clk, Q => 
                           n10728, QN => n8550);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2024, CK => Clk, Q => 
                           n10727, QN => n8551);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2023, CK => Clk, Q => n10726
                           , QN => n8552);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2022, CK => Clk, Q => n10725
                           , QN => n8553);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2021, CK => Clk, Q => n10724
                           , QN => n8554);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2020, CK => Clk, Q => n10723
                           , QN => n8555);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2019, CK => Clk, Q => n10722
                           , QN => n8556);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2018, CK => Clk, Q => n10721
                           , QN => n8557);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2017, CK => Clk, Q => n10720
                           , QN => n8558);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2016, CK => Clk, Q => n10719
                           , QN => n8559);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2015, CK => Clk, Q => n10718
                           , QN => n8560);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2014, CK => Clk, Q => n10717
                           , QN => n8561);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2069, CK => Clk, Q => 
                           n11124, QN => n8506);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2068, CK => Clk, Q => 
                           n11123, QN => n8507);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2067, CK => Clk, Q => 
                           n11122, QN => n8508);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2066, CK => Clk, Q => 
                           n11121, QN => n8509);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2065, CK => Clk, Q => 
                           n11120, QN => n8510);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2064, CK => Clk, Q => 
                           n11119, QN => n8511);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2063, CK => Clk, Q => 
                           n11118, QN => n8512);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2062, CK => Clk, Q => 
                           n11117, QN => n8513);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2061, CK => Clk, Q => 
                           n11116, QN => n8514);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2060, CK => Clk, Q => 
                           n11115, QN => n8515);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2059, CK => Clk, Q => 
                           n11114, QN => n8516);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2058, CK => Clk, Q => 
                           n11113, QN => n8517);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2057, CK => Clk, Q => 
                           n11112, QN => n8518);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2056, CK => Clk, Q => 
                           n11111, QN => n8519);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2055, CK => Clk, Q => n11110
                           , QN => n8520);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2054, CK => Clk, Q => n11109
                           , QN => n8521);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2053, CK => Clk, Q => n11108
                           , QN => n8522);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2052, CK => Clk, Q => n11107
                           , QN => n8523);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2051, CK => Clk, Q => n11106
                           , QN => n8524);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2050, CK => Clk, Q => n11105
                           , QN => n8525);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2049, CK => Clk, Q => n11104
                           , QN => n8526);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2048, CK => Clk, Q => n11103
                           , QN => n8527);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2047, CK => Clk, Q => n11102
                           , QN => n8528);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2046, CK => Clk, Q => n11101
                           , QN => n8529);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2197, CK => Clk, Q => 
                           n11188, QN => n8378);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2196, CK => Clk, Q => 
                           n11187, QN => n8379);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2195, CK => Clk, Q => 
                           n11186, QN => n8380);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2194, CK => Clk, Q => 
                           n11185, QN => n8381);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2193, CK => Clk, Q => 
                           n11184, QN => n8382);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2192, CK => Clk, Q => 
                           n11183, QN => n8383);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2191, CK => Clk, Q => 
                           n11182, QN => n8384);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2190, CK => Clk, Q => 
                           n11181, QN => n8385);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2189, CK => Clk, Q => 
                           n11180, QN => n8386);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2188, CK => Clk, Q => 
                           n11179, QN => n8387);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2187, CK => Clk, Q => 
                           n11178, QN => n8388);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2186, CK => Clk, Q => 
                           n11177, QN => n8389);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2185, CK => Clk, Q => 
                           n11176, QN => n8390);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2184, CK => Clk, Q => 
                           n11175, QN => n8391);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2183, CK => Clk, Q => n11174
                           , QN => n8392);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2182, CK => Clk, Q => n11173
                           , QN => n8393);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2181, CK => Clk, Q => n11172
                           , QN => n8394);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2180, CK => Clk, Q => n11171
                           , QN => n8395);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2179, CK => Clk, Q => n11170
                           , QN => n8396);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2178, CK => Clk, Q => n11169
                           , QN => n8397);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2177, CK => Clk, Q => n11168
                           , QN => n8398);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2176, CK => Clk, Q => n11167
                           , QN => n8399);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2175, CK => Clk, Q => n11166
                           , QN => n8400);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2174, CK => Clk, Q => n11165
                           , QN => n8401);
   Out2_reg_31_inst : DFF_X1 port map( D => n7245, CK => Clk, Q => Out2_31_port
                           , QN => n_1639);
   U7522 : BUF_X1 port map( A => n11419, Z => n11417);
   U7523 : BUF_X1 port map( A => n11607, Z => n11605);
   U7524 : BUF_X1 port map( A => n11419, Z => n11418);
   U7525 : BUF_X1 port map( A => n11607, Z => n11606);
   U7526 : BUF_X1 port map( A => n11359, Z => n11357);
   U7527 : BUF_X1 port map( A => n11363, Z => n11361);
   U7528 : BUF_X1 port map( A => n11367, Z => n11365);
   U7529 : BUF_X1 port map( A => n11371, Z => n11369);
   U7530 : BUF_X1 port map( A => n11375, Z => n11373);
   U7531 : BUF_X1 port map( A => n11379, Z => n11377);
   U7532 : BUF_X1 port map( A => n11383, Z => n11381);
   U7533 : BUF_X1 port map( A => n11387, Z => n11385);
   U7534 : BUF_X1 port map( A => n11391, Z => n11389);
   U7535 : BUF_X1 port map( A => n11395, Z => n11393);
   U7536 : BUF_X1 port map( A => n11399, Z => n11397);
   U7537 : BUF_X1 port map( A => n11403, Z => n11401);
   U7538 : BUF_X1 port map( A => n11407, Z => n11405);
   U7539 : BUF_X1 port map( A => n11411, Z => n11409);
   U7540 : BUF_X1 port map( A => n11415, Z => n11413);
   U7541 : BUF_X1 port map( A => n11423, Z => n11421);
   U7542 : BUF_X1 port map( A => n11427, Z => n11425);
   U7543 : BUF_X1 port map( A => n11431, Z => n11429);
   U7544 : BUF_X1 port map( A => n11435, Z => n11433);
   U7545 : BUF_X1 port map( A => n11439, Z => n11437);
   U7546 : BUF_X1 port map( A => n11443, Z => n11441);
   U7547 : BUF_X1 port map( A => n11447, Z => n11445);
   U7548 : BUF_X1 port map( A => n11451, Z => n11449);
   U7549 : BUF_X1 port map( A => n11455, Z => n11453);
   U7550 : BUF_X1 port map( A => n11459, Z => n11457);
   U7551 : BUF_X1 port map( A => n11463, Z => n11461);
   U7552 : BUF_X1 port map( A => n11467, Z => n11465);
   U7553 : BUF_X1 port map( A => n11471, Z => n11469);
   U7554 : BUF_X1 port map( A => n11475, Z => n11473);
   U7555 : BUF_X1 port map( A => n11479, Z => n11477);
   U7556 : BUF_X1 port map( A => n11359, Z => n11358);
   U7557 : BUF_X1 port map( A => n11363, Z => n11362);
   U7558 : BUF_X1 port map( A => n11367, Z => n11366);
   U7559 : BUF_X1 port map( A => n11371, Z => n11370);
   U7560 : BUF_X1 port map( A => n11375, Z => n11374);
   U7561 : BUF_X1 port map( A => n11379, Z => n11378);
   U7562 : BUF_X1 port map( A => n11383, Z => n11382);
   U7563 : BUF_X1 port map( A => n11387, Z => n11386);
   U7564 : BUF_X1 port map( A => n11391, Z => n11390);
   U7565 : BUF_X1 port map( A => n11395, Z => n11394);
   U7566 : BUF_X1 port map( A => n11399, Z => n11398);
   U7567 : BUF_X1 port map( A => n11403, Z => n11402);
   U7568 : BUF_X1 port map( A => n11407, Z => n11406);
   U7569 : BUF_X1 port map( A => n11411, Z => n11410);
   U7570 : BUF_X1 port map( A => n11415, Z => n11414);
   U7571 : BUF_X1 port map( A => n11423, Z => n11422);
   U7572 : BUF_X1 port map( A => n11427, Z => n11426);
   U7573 : BUF_X1 port map( A => n11431, Z => n11430);
   U7574 : BUF_X1 port map( A => n11435, Z => n11434);
   U7575 : BUF_X1 port map( A => n11439, Z => n11438);
   U7576 : BUF_X1 port map( A => n11443, Z => n11442);
   U7577 : BUF_X1 port map( A => n11447, Z => n11446);
   U7578 : BUF_X1 port map( A => n11451, Z => n11450);
   U7579 : BUF_X1 port map( A => n11455, Z => n11454);
   U7580 : BUF_X1 port map( A => n11459, Z => n11458);
   U7581 : BUF_X1 port map( A => n11463, Z => n11462);
   U7582 : BUF_X1 port map( A => n11467, Z => n11466);
   U7583 : BUF_X1 port map( A => n11471, Z => n11470);
   U7584 : BUF_X1 port map( A => n11475, Z => n11474);
   U7585 : BUF_X1 port map( A => n11479, Z => n11478);
   U7586 : BUF_X1 port map( A => n9895, Z => n11742);
   U7587 : BUF_X1 port map( A => n9305, Z => n11881);
   U7588 : BUF_X1 port map( A => n9896, Z => n11738);
   U7589 : BUF_X1 port map( A => n9306, Z => n11877);
   U7590 : BUF_X1 port map( A => n9900, Z => n11726);
   U7591 : BUF_X1 port map( A => n9906, Z => n11706);
   U7592 : BUF_X1 port map( A => n9310, Z => n11865);
   U7593 : BUF_X1 port map( A => n9316, Z => n11845);
   U7594 : BUF_X1 port map( A => n9911, Z => n11691);
   U7595 : BUF_X1 port map( A => n9905, Z => n11710);
   U7596 : BUF_X1 port map( A => n9321, Z => n11830);
   U7597 : BUF_X1 port map( A => n9315, Z => n11849);
   U7598 : BUF_X1 port map( A => n9912, Z => n11687);
   U7599 : BUF_X1 port map( A => n9901, Z => n11722);
   U7600 : BUF_X1 port map( A => n9322, Z => n11826);
   U7601 : BUF_X1 port map( A => n9311, Z => n11861);
   U7602 : BUF_X1 port map( A => n8260, Z => n11896);
   U7603 : BUF_X1 port map( A => n8260, Z => n11897);
   U7604 : BUF_X1 port map( A => n9892, Z => n11747);
   U7605 : BUF_X1 port map( A => n9893, Z => n11743);
   U7606 : BUF_X1 port map( A => n9897, Z => n11731);
   U7607 : BUF_X1 port map( A => n9898, Z => n11727);
   U7608 : BUF_X1 port map( A => n9902, Z => n11715);
   U7609 : BUF_X1 port map( A => n9903, Z => n11711);
   U7610 : BUF_X1 port map( A => n9303, Z => n11882);
   U7611 : BUF_X1 port map( A => n9302, Z => n11886);
   U7612 : BUF_X1 port map( A => n9308, Z => n11866);
   U7613 : BUF_X1 port map( A => n9307, Z => n11870);
   U7614 : BUF_X1 port map( A => n9313, Z => n11850);
   U7615 : BUF_X1 port map( A => n9312, Z => n11854);
   U7616 : BUF_X1 port map( A => n9921, Z => n11668);
   U7617 : BUF_X1 port map( A => n9937, Z => n11616);
   U7618 : BUF_X1 port map( A => n9938, Z => n11612);
   U7619 : BUF_X1 port map( A => n11702, Z => n11700);
   U7620 : BUF_X1 port map( A => n9331, Z => n11807);
   U7621 : BUF_X1 port map( A => n9348, Z => n11751);
   U7622 : BUF_X1 port map( A => n9347, Z => n11755);
   U7623 : BUF_X1 port map( A => n11841, Z => n11839);
   U7624 : BUF_X1 port map( A => n9917, Z => n11680);
   U7625 : BUF_X1 port map( A => n9918, Z => n11676);
   U7626 : BUF_X1 port map( A => n9928, Z => n11644);
   U7627 : BUF_X1 port map( A => n9929, Z => n11640);
   U7628 : BUF_X1 port map( A => n9923, Z => n11660);
   U7629 : BUF_X1 port map( A => n9924, Z => n11656);
   U7630 : BUF_X1 port map( A => n9934, Z => n11624);
   U7631 : BUF_X1 port map( A => n9935, Z => n11620);
   U7632 : BUF_X1 port map( A => n9328, Z => n11815);
   U7633 : BUF_X1 port map( A => n9327, Z => n11819);
   U7634 : BUF_X1 port map( A => n9339, Z => n11779);
   U7635 : BUF_X1 port map( A => n9338, Z => n11783);
   U7636 : BUF_X1 port map( A => n9334, Z => n11795);
   U7637 : BUF_X1 port map( A => n9333, Z => n11799);
   U7638 : BUF_X1 port map( A => n9345, Z => n11759);
   U7639 : BUF_X1 port map( A => n9344, Z => n11763);
   U7640 : BUF_X1 port map( A => n9922, Z => n11664);
   U7641 : BUF_X1 port map( A => n9920, Z => n11672);
   U7642 : BUF_X1 port map( A => n9933, Z => n11628);
   U7643 : BUF_X1 port map( A => n9932, Z => n11632);
   U7644 : BUF_X1 port map( A => n9931, Z => n11636);
   U7645 : BUF_X1 port map( A => n9926, Z => n11652);
   U7646 : BUF_X1 port map( A => n9927, Z => n11648);
   U7647 : BUF_X1 port map( A => n9332, Z => n11803);
   U7648 : BUF_X1 port map( A => n9330, Z => n11811);
   U7649 : BUF_X1 port map( A => n9343, Z => n11767);
   U7650 : BUF_X1 port map( A => n9342, Z => n11771);
   U7651 : BUF_X1 port map( A => n9341, Z => n11775);
   U7652 : BUF_X1 port map( A => n9337, Z => n11787);
   U7653 : BUF_X1 port map( A => n9336, Z => n11791);
   U7654 : BUF_X1 port map( A => n9909, Z => n11695);
   U7655 : BUF_X1 port map( A => n9319, Z => n11834);
   U7656 : BUF_X1 port map( A => n10510, Z => n11480);
   U7657 : BUF_X1 port map( A => n10509, Z => n11484);
   U7658 : BUF_X1 port map( A => n10508, Z => n11488);
   U7659 : BUF_X1 port map( A => n10507, Z => n11492);
   U7660 : BUF_X1 port map( A => n10506, Z => n11496);
   U7661 : BUF_X1 port map( A => n10505, Z => n11500);
   U7662 : BUF_X1 port map( A => n10504, Z => n11504);
   U7663 : BUF_X1 port map( A => n10503, Z => n11508);
   U7664 : BUF_X1 port map( A => n10502, Z => n11512);
   U7665 : BUF_X1 port map( A => n10501, Z => n11516);
   U7666 : BUF_X1 port map( A => n10500, Z => n11520);
   U7667 : BUF_X1 port map( A => n10499, Z => n11524);
   U7668 : BUF_X1 port map( A => n10498, Z => n11528);
   U7669 : BUF_X1 port map( A => n10497, Z => n11532);
   U7670 : BUF_X1 port map( A => n10496, Z => n11536);
   U7671 : BUF_X1 port map( A => n10495, Z => n11540);
   U7672 : BUF_X1 port map( A => n10494, Z => n11544);
   U7673 : BUF_X1 port map( A => n10493, Z => n11548);
   U7674 : BUF_X1 port map( A => n10492, Z => n11552);
   U7675 : BUF_X1 port map( A => n10491, Z => n11556);
   U7676 : BUF_X1 port map( A => n10490, Z => n11560);
   U7677 : BUF_X1 port map( A => n10489, Z => n11564);
   U7678 : BUF_X1 port map( A => n10488, Z => n11568);
   U7679 : BUF_X1 port map( A => n10487, Z => n11572);
   U7680 : BUF_X1 port map( A => n10486, Z => n11576);
   U7681 : BUF_X1 port map( A => n10485, Z => n11580);
   U7682 : BUF_X1 port map( A => n10484, Z => n11584);
   U7683 : BUF_X1 port map( A => n10483, Z => n11588);
   U7684 : BUF_X1 port map( A => n10482, Z => n11592);
   U7685 : BUF_X1 port map( A => n10481, Z => n11596);
   U7686 : BUF_X1 port map( A => n10480, Z => n11600);
   U7687 : BUF_X1 port map( A => n10478, Z => n11608);
   U7688 : BUF_X1 port map( A => n11418, Z => n11306);
   U7689 : BUF_X1 port map( A => n11418, Z => n11305);
   U7690 : BUF_X1 port map( A => n11606, Z => n11354);
   U7691 : BUF_X1 port map( A => n11606, Z => n11353);
   U7692 : INV_X1 port map( A => n11417, ZN => n11416);
   U7693 : INV_X1 port map( A => n11605, ZN => n11604);
   U7694 : BUF_X1 port map( A => n11418, Z => n11307);
   U7695 : BUF_X1 port map( A => n11606, Z => n11355);
   U7696 : BUF_X1 port map( A => n11358, Z => n11261);
   U7697 : BUF_X1 port map( A => n11358, Z => n11260);
   U7698 : BUF_X1 port map( A => n11362, Z => n11264);
   U7699 : BUF_X1 port map( A => n11362, Z => n11263);
   U7700 : BUF_X1 port map( A => n11366, Z => n11267);
   U7701 : BUF_X1 port map( A => n11366, Z => n11266);
   U7702 : BUF_X1 port map( A => n11370, Z => n11270);
   U7703 : BUF_X1 port map( A => n11370, Z => n11269);
   U7704 : BUF_X1 port map( A => n11374, Z => n11273);
   U7705 : BUF_X1 port map( A => n11374, Z => n11272);
   U7706 : BUF_X1 port map( A => n11378, Z => n11276);
   U7707 : BUF_X1 port map( A => n11378, Z => n11275);
   U7708 : BUF_X1 port map( A => n11382, Z => n11279);
   U7709 : BUF_X1 port map( A => n11382, Z => n11278);
   U7710 : BUF_X1 port map( A => n11386, Z => n11282);
   U7711 : BUF_X1 port map( A => n11386, Z => n11281);
   U7712 : BUF_X1 port map( A => n11390, Z => n11285);
   U7713 : BUF_X1 port map( A => n11390, Z => n11284);
   U7714 : BUF_X1 port map( A => n11394, Z => n11288);
   U7715 : BUF_X1 port map( A => n11394, Z => n11287);
   U7716 : BUF_X1 port map( A => n11398, Z => n11291);
   U7717 : BUF_X1 port map( A => n11398, Z => n11290);
   U7718 : BUF_X1 port map( A => n11402, Z => n11294);
   U7719 : BUF_X1 port map( A => n11402, Z => n11293);
   U7720 : BUF_X1 port map( A => n11406, Z => n11297);
   U7721 : BUF_X1 port map( A => n11406, Z => n11296);
   U7722 : BUF_X1 port map( A => n11410, Z => n11300);
   U7723 : BUF_X1 port map( A => n11410, Z => n11299);
   U7724 : BUF_X1 port map( A => n11414, Z => n11303);
   U7725 : BUF_X1 port map( A => n11414, Z => n11302);
   U7726 : BUF_X1 port map( A => n11422, Z => n11309);
   U7727 : BUF_X1 port map( A => n11422, Z => n11308);
   U7728 : BUF_X1 port map( A => n11426, Z => n11312);
   U7729 : BUF_X1 port map( A => n11426, Z => n11311);
   U7730 : BUF_X1 port map( A => n11430, Z => n11315);
   U7731 : BUF_X1 port map( A => n11430, Z => n11314);
   U7732 : BUF_X1 port map( A => n11434, Z => n11318);
   U7733 : BUF_X1 port map( A => n11434, Z => n11317);
   U7734 : BUF_X1 port map( A => n11438, Z => n11321);
   U7735 : BUF_X1 port map( A => n11438, Z => n11320);
   U7736 : BUF_X1 port map( A => n11442, Z => n11324);
   U7737 : BUF_X1 port map( A => n11442, Z => n11323);
   U7738 : BUF_X1 port map( A => n11446, Z => n11327);
   U7739 : BUF_X1 port map( A => n11446, Z => n11326);
   U7740 : BUF_X1 port map( A => n11450, Z => n11330);
   U7741 : BUF_X1 port map( A => n11450, Z => n11329);
   U7742 : BUF_X1 port map( A => n11454, Z => n11333);
   U7743 : BUF_X1 port map( A => n11454, Z => n11332);
   U7744 : BUF_X1 port map( A => n11458, Z => n11336);
   U7745 : BUF_X1 port map( A => n11458, Z => n11335);
   U7746 : BUF_X1 port map( A => n11462, Z => n11339);
   U7747 : BUF_X1 port map( A => n11462, Z => n11338);
   U7748 : BUF_X1 port map( A => n11466, Z => n11342);
   U7749 : BUF_X1 port map( A => n11466, Z => n11341);
   U7750 : BUF_X1 port map( A => n11470, Z => n11345);
   U7751 : BUF_X1 port map( A => n11470, Z => n11344);
   U7752 : BUF_X1 port map( A => n11474, Z => n11348);
   U7753 : BUF_X1 port map( A => n11474, Z => n11347);
   U7754 : BUF_X1 port map( A => n11478, Z => n11351);
   U7755 : BUF_X1 port map( A => n11478, Z => n11350);
   U7756 : INV_X1 port map( A => n11357, ZN => n11356);
   U7757 : INV_X1 port map( A => n11361, ZN => n11360);
   U7758 : INV_X1 port map( A => n11365, ZN => n11364);
   U7759 : INV_X1 port map( A => n11369, ZN => n11368);
   U7760 : INV_X1 port map( A => n11373, ZN => n11372);
   U7761 : INV_X1 port map( A => n11377, ZN => n11376);
   U7762 : INV_X1 port map( A => n11381, ZN => n11380);
   U7763 : INV_X1 port map( A => n11385, ZN => n11384);
   U7764 : INV_X1 port map( A => n11389, ZN => n11388);
   U7765 : INV_X1 port map( A => n11393, ZN => n11392);
   U7766 : INV_X1 port map( A => n11397, ZN => n11396);
   U7767 : INV_X1 port map( A => n11401, ZN => n11400);
   U7768 : INV_X1 port map( A => n11405, ZN => n11404);
   U7769 : INV_X1 port map( A => n11409, ZN => n11408);
   U7770 : INV_X1 port map( A => n11413, ZN => n11412);
   U7771 : INV_X1 port map( A => n11421, ZN => n11420);
   U7772 : INV_X1 port map( A => n11425, ZN => n11424);
   U7773 : INV_X1 port map( A => n11429, ZN => n11428);
   U7774 : INV_X1 port map( A => n11433, ZN => n11432);
   U7775 : INV_X1 port map( A => n11437, ZN => n11436);
   U7776 : INV_X1 port map( A => n11441, ZN => n11440);
   U7777 : INV_X1 port map( A => n11445, ZN => n11444);
   U7778 : INV_X1 port map( A => n11449, ZN => n11448);
   U7779 : INV_X1 port map( A => n11453, ZN => n11452);
   U7780 : INV_X1 port map( A => n11457, ZN => n11456);
   U7781 : INV_X1 port map( A => n11461, ZN => n11460);
   U7782 : INV_X1 port map( A => n11465, ZN => n11464);
   U7783 : INV_X1 port map( A => n11469, ZN => n11468);
   U7784 : INV_X1 port map( A => n11473, ZN => n11472);
   U7785 : INV_X1 port map( A => n11477, ZN => n11476);
   U7786 : BUF_X1 port map( A => n11358, Z => n11262);
   U7787 : BUF_X1 port map( A => n11362, Z => n11265);
   U7788 : BUF_X1 port map( A => n11366, Z => n11268);
   U7789 : BUF_X1 port map( A => n11370, Z => n11271);
   U7790 : BUF_X1 port map( A => n11374, Z => n11274);
   U7791 : BUF_X1 port map( A => n11378, Z => n11277);
   U7792 : BUF_X1 port map( A => n11382, Z => n11280);
   U7793 : BUF_X1 port map( A => n11386, Z => n11283);
   U7794 : BUF_X1 port map( A => n11390, Z => n11286);
   U7795 : BUF_X1 port map( A => n11394, Z => n11289);
   U7796 : BUF_X1 port map( A => n11398, Z => n11292);
   U7797 : BUF_X1 port map( A => n11402, Z => n11295);
   U7798 : BUF_X1 port map( A => n11406, Z => n11298);
   U7799 : BUF_X1 port map( A => n11410, Z => n11301);
   U7800 : BUF_X1 port map( A => n11414, Z => n11304);
   U7801 : BUF_X1 port map( A => n11422, Z => n11310);
   U7802 : BUF_X1 port map( A => n11426, Z => n11313);
   U7803 : BUF_X1 port map( A => n11430, Z => n11316);
   U7804 : BUF_X1 port map( A => n11434, Z => n11319);
   U7805 : BUF_X1 port map( A => n11438, Z => n11322);
   U7806 : BUF_X1 port map( A => n11442, Z => n11325);
   U7807 : BUF_X1 port map( A => n11446, Z => n11328);
   U7808 : BUF_X1 port map( A => n11450, Z => n11331);
   U7809 : BUF_X1 port map( A => n11454, Z => n11334);
   U7810 : BUF_X1 port map( A => n11458, Z => n11337);
   U7811 : BUF_X1 port map( A => n11462, Z => n11340);
   U7812 : BUF_X1 port map( A => n11466, Z => n11343);
   U7813 : BUF_X1 port map( A => n11470, Z => n11346);
   U7814 : BUF_X1 port map( A => n11474, Z => n11349);
   U7815 : BUF_X1 port map( A => n11478, Z => n11352);
   U7816 : INV_X1 port map( A => n10535, ZN => n11419);
   U7817 : OAI21_X1 port map( B1 => n10512, B2 => n10536, A => n11893, ZN => 
                           n10535);
   U7818 : INV_X1 port map( A => n10479, ZN => n11607);
   U7819 : OAI21_X1 port map( B1 => n10511, B2 => n10512, A => n11892, ZN => 
                           n10479);
   U7820 : BUF_X1 port map( A => n11896, Z => n11893);
   U7821 : BUF_X1 port map( A => n11896, Z => n11894);
   U7822 : BUF_X1 port map( A => n11815, Z => n11816);
   U7823 : BUF_X1 port map( A => n11779, Z => n11780);
   U7824 : BUF_X1 port map( A => n11795, Z => n11796);
   U7825 : BUF_X1 port map( A => n11759, Z => n11760);
   U7826 : BUF_X1 port map( A => n11815, Z => n11817);
   U7827 : BUF_X1 port map( A => n11779, Z => n11781);
   U7828 : BUF_X1 port map( A => n11795, Z => n11797);
   U7829 : BUF_X1 port map( A => n11759, Z => n11761);
   U7830 : BUF_X1 port map( A => n11882, Z => n11883);
   U7831 : BUF_X1 port map( A => n11866, Z => n11867);
   U7832 : BUF_X1 port map( A => n11850, Z => n11851);
   U7833 : BUF_X1 port map( A => n11882, Z => n11884);
   U7834 : BUF_X1 port map( A => n11866, Z => n11868);
   U7835 : BUF_X1 port map( A => n11850, Z => n11852);
   U7836 : BUF_X1 port map( A => n11897, Z => n11891);
   U7837 : BUF_X1 port map( A => n11897, Z => n11890);
   U7838 : BUF_X1 port map( A => n11691, Z => n11688);
   U7839 : BUF_X1 port map( A => n11742, Z => n11739);
   U7840 : BUF_X1 port map( A => n11726, Z => n11723);
   U7841 : BUF_X1 port map( A => n11710, Z => n11707);
   U7842 : BUF_X1 port map( A => n11691, Z => n11689);
   U7843 : BUF_X1 port map( A => n11742, Z => n11740);
   U7844 : BUF_X1 port map( A => n11726, Z => n11724);
   U7845 : BUF_X1 port map( A => n11710, Z => n11708);
   U7846 : BUF_X1 port map( A => n11652, Z => n11653);
   U7847 : BUF_X1 port map( A => n11616, Z => n11617);
   U7848 : BUF_X1 port map( A => n11652, Z => n11654);
   U7849 : BUF_X1 port map( A => n11616, Z => n11618);
   U7850 : BUF_X1 port map( A => n11803, Z => n11804);
   U7851 : BUF_X1 port map( A => n11767, Z => n11768);
   U7852 : BUF_X1 port map( A => n11803, Z => n11805);
   U7853 : BUF_X1 port map( A => n11767, Z => n11769);
   U7854 : BUF_X1 port map( A => n11897, Z => n11892);
   U7855 : BUF_X1 port map( A => n11687, Z => n11684);
   U7856 : BUF_X1 port map( A => n11738, Z => n11735);
   U7857 : BUF_X1 port map( A => n11722, Z => n11719);
   U7858 : BUF_X1 port map( A => n11706, Z => n11703);
   U7859 : BUF_X1 port map( A => n11687, Z => n11685);
   U7860 : BUF_X1 port map( A => n11738, Z => n11736);
   U7861 : BUF_X1 port map( A => n11722, Z => n11720);
   U7862 : BUF_X1 port map( A => n11706, Z => n11704);
   U7863 : BUF_X1 port map( A => n11648, Z => n11649);
   U7864 : BUF_X1 port map( A => n11612, Z => n11613);
   U7865 : BUF_X1 port map( A => n11648, Z => n11650);
   U7866 : BUF_X1 port map( A => n11612, Z => n11614);
   U7867 : BUF_X1 port map( A => n11807, Z => n11808);
   U7868 : BUF_X1 port map( A => n11771, Z => n11772);
   U7869 : BUF_X1 port map( A => n11807, Z => n11809);
   U7870 : BUF_X1 port map( A => n11771, Z => n11773);
   U7871 : BUF_X1 port map( A => n11811, Z => n11812);
   U7872 : BUF_X1 port map( A => n11775, Z => n11776);
   U7873 : BUF_X1 port map( A => n11811, Z => n11813);
   U7874 : BUF_X1 port map( A => n11775, Z => n11777);
   U7875 : BUF_X1 port map( A => n11680, Z => n11681);
   U7876 : BUF_X1 port map( A => n11644, Z => n11645);
   U7877 : BUF_X1 port map( A => n11660, Z => n11661);
   U7878 : BUF_X1 port map( A => n11624, Z => n11625);
   U7879 : BUF_X1 port map( A => n11680, Z => n11682);
   U7880 : BUF_X1 port map( A => n11644, Z => n11646);
   U7881 : BUF_X1 port map( A => n11660, Z => n11662);
   U7882 : BUF_X1 port map( A => n11624, Z => n11626);
   U7883 : BUF_X1 port map( A => n11747, Z => n11748);
   U7884 : BUF_X1 port map( A => n11731, Z => n11732);
   U7885 : BUF_X1 port map( A => n11715, Z => n11716);
   U7886 : BUF_X1 port map( A => n11747, Z => n11749);
   U7887 : BUF_X1 port map( A => n11731, Z => n11733);
   U7888 : BUF_X1 port map( A => n11715, Z => n11717);
   U7889 : BUF_X1 port map( A => n11700, Z => n11697);
   U7890 : BUF_X1 port map( A => n11839, Z => n11836);
   U7891 : BUF_X1 port map( A => n11826, Z => n11823);
   U7892 : BUF_X1 port map( A => n11877, Z => n11874);
   U7893 : BUF_X1 port map( A => n11861, Z => n11858);
   U7894 : BUF_X1 port map( A => n11845, Z => n11842);
   U7895 : BUF_X1 port map( A => n11826, Z => n11824);
   U7896 : BUF_X1 port map( A => n11877, Z => n11875);
   U7897 : BUF_X1 port map( A => n11861, Z => n11859);
   U7898 : BUF_X1 port map( A => n11845, Z => n11843);
   U7899 : BUF_X1 port map( A => n11787, Z => n11788);
   U7900 : BUF_X1 port map( A => n11751, Z => n11752);
   U7901 : BUF_X1 port map( A => n11787, Z => n11789);
   U7902 : BUF_X1 port map( A => n11751, Z => n11753);
   U7903 : BUF_X1 port map( A => n11830, Z => n11827);
   U7904 : BUF_X1 port map( A => n11881, Z => n11878);
   U7905 : BUF_X1 port map( A => n11865, Z => n11862);
   U7906 : BUF_X1 port map( A => n11849, Z => n11846);
   U7907 : BUF_X1 port map( A => n11830, Z => n11828);
   U7908 : BUF_X1 port map( A => n11881, Z => n11879);
   U7909 : BUF_X1 port map( A => n11865, Z => n11863);
   U7910 : BUF_X1 port map( A => n11849, Z => n11847);
   U7911 : BUF_X1 port map( A => n11676, Z => n11677);
   U7912 : BUF_X1 port map( A => n11640, Z => n11641);
   U7913 : BUF_X1 port map( A => n11656, Z => n11657);
   U7914 : BUF_X1 port map( A => n11620, Z => n11621);
   U7915 : BUF_X1 port map( A => n11676, Z => n11678);
   U7916 : BUF_X1 port map( A => n11640, Z => n11642);
   U7917 : BUF_X1 port map( A => n11656, Z => n11658);
   U7918 : BUF_X1 port map( A => n11620, Z => n11622);
   U7919 : BUF_X1 port map( A => n11743, Z => n11744);
   U7920 : BUF_X1 port map( A => n11727, Z => n11728);
   U7921 : BUF_X1 port map( A => n11711, Z => n11712);
   U7922 : BUF_X1 port map( A => n11743, Z => n11745);
   U7923 : BUF_X1 port map( A => n11727, Z => n11729);
   U7924 : BUF_X1 port map( A => n11711, Z => n11713);
   U7925 : BUF_X1 port map( A => n11819, Z => n11820);
   U7926 : BUF_X1 port map( A => n11783, Z => n11784);
   U7927 : BUF_X1 port map( A => n11799, Z => n11800);
   U7928 : BUF_X1 port map( A => n11763, Z => n11764);
   U7929 : BUF_X1 port map( A => n11819, Z => n11821);
   U7930 : BUF_X1 port map( A => n11783, Z => n11785);
   U7931 : BUF_X1 port map( A => n11799, Z => n11801);
   U7932 : BUF_X1 port map( A => n11763, Z => n11765);
   U7933 : BUF_X1 port map( A => n11886, Z => n11887);
   U7934 : BUF_X1 port map( A => n11870, Z => n11871);
   U7935 : BUF_X1 port map( A => n11854, Z => n11855);
   U7936 : BUF_X1 port map( A => n11886, Z => n11888);
   U7937 : BUF_X1 port map( A => n11870, Z => n11872);
   U7938 : BUF_X1 port map( A => n11854, Z => n11856);
   U7939 : BUF_X1 port map( A => n11791, Z => n11792);
   U7940 : BUF_X1 port map( A => n11755, Z => n11756);
   U7941 : BUF_X1 port map( A => n11791, Z => n11793);
   U7942 : BUF_X1 port map( A => n11755, Z => n11757);
   U7943 : BUF_X1 port map( A => n11700, Z => n11698);
   U7944 : BUF_X1 port map( A => n11839, Z => n11837);
   U7945 : BUF_X1 port map( A => n11664, Z => n11665);
   U7946 : BUF_X1 port map( A => n11628, Z => n11629);
   U7947 : BUF_X1 port map( A => n11664, Z => n11666);
   U7948 : BUF_X1 port map( A => n11628, Z => n11630);
   U7949 : BUF_X1 port map( A => n11668, Z => n11669);
   U7950 : BUF_X1 port map( A => n11632, Z => n11633);
   U7951 : BUF_X1 port map( A => n11668, Z => n11670);
   U7952 : BUF_X1 port map( A => n11632, Z => n11634);
   U7953 : BUF_X1 port map( A => n11672, Z => n11673);
   U7954 : BUF_X1 port map( A => n11636, Z => n11637);
   U7955 : BUF_X1 port map( A => n11672, Z => n11674);
   U7956 : BUF_X1 port map( A => n11636, Z => n11638);
   U7957 : BUF_X1 port map( A => n11815, Z => n11818);
   U7958 : BUF_X1 port map( A => n11779, Z => n11782);
   U7959 : BUF_X1 port map( A => n11795, Z => n11798);
   U7960 : BUF_X1 port map( A => n11759, Z => n11762);
   U7961 : BUF_X1 port map( A => n11882, Z => n11885);
   U7962 : BUF_X1 port map( A => n11866, Z => n11869);
   U7963 : BUF_X1 port map( A => n11850, Z => n11853);
   U7964 : BUF_X1 port map( A => n11691, Z => n11690);
   U7965 : BUF_X1 port map( A => n11742, Z => n11741);
   U7966 : BUF_X1 port map( A => n11726, Z => n11725);
   U7967 : BUF_X1 port map( A => n11710, Z => n11709);
   U7968 : BUF_X1 port map( A => n11652, Z => n11655);
   U7969 : BUF_X1 port map( A => n11616, Z => n11619);
   U7970 : BUF_X1 port map( A => n11803, Z => n11806);
   U7971 : BUF_X1 port map( A => n11767, Z => n11770);
   U7972 : BUF_X1 port map( A => n11687, Z => n11686);
   U7973 : BUF_X1 port map( A => n11738, Z => n11737);
   U7974 : BUF_X1 port map( A => n11722, Z => n11721);
   U7975 : BUF_X1 port map( A => n11706, Z => n11705);
   U7976 : BUF_X1 port map( A => n11648, Z => n11651);
   U7977 : BUF_X1 port map( A => n11612, Z => n11615);
   U7978 : BUF_X1 port map( A => n11807, Z => n11810);
   U7979 : BUF_X1 port map( A => n11771, Z => n11774);
   U7980 : BUF_X1 port map( A => n11811, Z => n11814);
   U7981 : BUF_X1 port map( A => n11775, Z => n11778);
   U7982 : BUF_X1 port map( A => n11680, Z => n11683);
   U7983 : BUF_X1 port map( A => n11644, Z => n11647);
   U7984 : BUF_X1 port map( A => n11660, Z => n11663);
   U7985 : BUF_X1 port map( A => n11624, Z => n11627);
   U7986 : BUF_X1 port map( A => n11747, Z => n11750);
   U7987 : BUF_X1 port map( A => n11731, Z => n11734);
   U7988 : BUF_X1 port map( A => n11715, Z => n11718);
   U7989 : BUF_X1 port map( A => n11826, Z => n11825);
   U7990 : BUF_X1 port map( A => n11877, Z => n11876);
   U7991 : BUF_X1 port map( A => n11861, Z => n11860);
   U7992 : BUF_X1 port map( A => n11845, Z => n11844);
   U7993 : BUF_X1 port map( A => n11830, Z => n11829);
   U7994 : BUF_X1 port map( A => n11881, Z => n11880);
   U7995 : BUF_X1 port map( A => n11865, Z => n11864);
   U7996 : BUF_X1 port map( A => n11849, Z => n11848);
   U7997 : BUF_X1 port map( A => n11787, Z => n11790);
   U7998 : BUF_X1 port map( A => n11751, Z => n11754);
   U7999 : BUF_X1 port map( A => n11676, Z => n11679);
   U8000 : BUF_X1 port map( A => n11640, Z => n11643);
   U8001 : BUF_X1 port map( A => n11656, Z => n11659);
   U8002 : BUF_X1 port map( A => n11620, Z => n11623);
   U8003 : BUF_X1 port map( A => n11743, Z => n11746);
   U8004 : BUF_X1 port map( A => n11727, Z => n11730);
   U8005 : BUF_X1 port map( A => n11711, Z => n11714);
   U8006 : BUF_X1 port map( A => n11819, Z => n11822);
   U8007 : BUF_X1 port map( A => n11783, Z => n11786);
   U8008 : BUF_X1 port map( A => n11799, Z => n11802);
   U8009 : BUF_X1 port map( A => n11763, Z => n11766);
   U8010 : BUF_X1 port map( A => n11886, Z => n11889);
   U8011 : BUF_X1 port map( A => n11870, Z => n11873);
   U8012 : BUF_X1 port map( A => n11854, Z => n11857);
   U8013 : BUF_X1 port map( A => n11791, Z => n11794);
   U8014 : BUF_X1 port map( A => n11755, Z => n11758);
   U8015 : BUF_X1 port map( A => n11664, Z => n11667);
   U8016 : BUF_X1 port map( A => n11628, Z => n11631);
   U8017 : BUF_X1 port map( A => n11668, Z => n11671);
   U8018 : BUF_X1 port map( A => n11632, Z => n11635);
   U8019 : BUF_X1 port map( A => n11672, Z => n11675);
   U8020 : BUF_X1 port map( A => n11636, Z => n11639);
   U8021 : BUF_X1 port map( A => n11700, Z => n11699);
   U8022 : BUF_X1 port map( A => n11839, Z => n11838);
   U8023 : BUF_X1 port map( A => n11896, Z => n11895);
   U8024 : OAI22_X1 port map( A1 => n11756, A2 => n9233, B1 => n11752, B2 => 
                           n8977, ZN => n9887);
   U8025 : OAI22_X1 port map( A1 => n11756, A2 => n9232, B1 => n11752, B2 => 
                           n8976, ZN => n9858);
   U8026 : OAI22_X1 port map( A1 => n11756, A2 => n9231, B1 => n11752, B2 => 
                           n8975, ZN => n9841);
   U8027 : OAI22_X1 port map( A1 => n11756, A2 => n9230, B1 => n11752, B2 => 
                           n8974, ZN => n9824);
   U8028 : OAI22_X1 port map( A1 => n11756, A2 => n9229, B1 => n11752, B2 => 
                           n8973, ZN => n9807);
   U8029 : OAI22_X1 port map( A1 => n11756, A2 => n9228, B1 => n11752, B2 => 
                           n8972, ZN => n9790);
   U8030 : OAI22_X1 port map( A1 => n11756, A2 => n9227, B1 => n11752, B2 => 
                           n8971, ZN => n9773);
   U8031 : OAI22_X1 port map( A1 => n11756, A2 => n9226, B1 => n11752, B2 => 
                           n8970, ZN => n9756);
   U8032 : OAI22_X1 port map( A1 => n11756, A2 => n9225, B1 => n11752, B2 => 
                           n8969, ZN => n9739);
   U8033 : OAI22_X1 port map( A1 => n11756, A2 => n9224, B1 => n11752, B2 => 
                           n8968, ZN => n9722);
   U8034 : OAI22_X1 port map( A1 => n11756, A2 => n9223, B1 => n11752, B2 => 
                           n8967, ZN => n9705);
   U8035 : OAI22_X1 port map( A1 => n11756, A2 => n9222, B1 => n11752, B2 => 
                           n8966, ZN => n9688);
   U8036 : OAI22_X1 port map( A1 => n11757, A2 => n9221, B1 => n11753, B2 => 
                           n8965, ZN => n9671);
   U8037 : OAI22_X1 port map( A1 => n11757, A2 => n9220, B1 => n11753, B2 => 
                           n8964, ZN => n9654);
   U8038 : OAI22_X1 port map( A1 => n11757, A2 => n9219, B1 => n11753, B2 => 
                           n8963, ZN => n9637);
   U8039 : OAI22_X1 port map( A1 => n11757, A2 => n9218, B1 => n11753, B2 => 
                           n8962, ZN => n9620);
   U8040 : OAI22_X1 port map( A1 => n11757, A2 => n9217, B1 => n11753, B2 => 
                           n8961, ZN => n9603);
   U8041 : OAI22_X1 port map( A1 => n11757, A2 => n9216, B1 => n11753, B2 => 
                           n8960, ZN => n9586);
   U8042 : OAI22_X1 port map( A1 => n11757, A2 => n9215, B1 => n11753, B2 => 
                           n8959, ZN => n9569);
   U8043 : OAI22_X1 port map( A1 => n11757, A2 => n9214, B1 => n11753, B2 => 
                           n8958, ZN => n9552);
   U8044 : OAI22_X1 port map( A1 => n11757, A2 => n9213, B1 => n11753, B2 => 
                           n8957, ZN => n9535);
   U8045 : OAI22_X1 port map( A1 => n11757, A2 => n9212, B1 => n11753, B2 => 
                           n8956, ZN => n9518);
   U8046 : OAI22_X1 port map( A1 => n11757, A2 => n9211, B1 => n11753, B2 => 
                           n8955, ZN => n9501);
   U8047 : OAI22_X1 port map( A1 => n11757, A2 => n9210, B1 => n11753, B2 => 
                           n8954, ZN => n9484);
   U8048 : OAI22_X1 port map( A1 => n11758, A2 => n9209, B1 => n11754, B2 => 
                           n8953, ZN => n9467);
   U8049 : OAI22_X1 port map( A1 => n11758, A2 => n9208, B1 => n11754, B2 => 
                           n8952, ZN => n9450);
   U8050 : OAI22_X1 port map( A1 => n11758, A2 => n9207, B1 => n11754, B2 => 
                           n8951, ZN => n9433);
   U8051 : OAI22_X1 port map( A1 => n11758, A2 => n9206, B1 => n11754, B2 => 
                           n8950, ZN => n9416);
   U8052 : OAI22_X1 port map( A1 => n11758, A2 => n9205, B1 => n11754, B2 => 
                           n8949, ZN => n9399);
   U8053 : OAI22_X1 port map( A1 => n11758, A2 => n9204, B1 => n11754, B2 => 
                           n8948, ZN => n9382);
   U8054 : OAI22_X1 port map( A1 => n11758, A2 => n9203, B1 => n11754, B2 => 
                           n8947, ZN => n9365);
   U8055 : OAI22_X1 port map( A1 => n11758, A2 => n9202, B1 => n11754, B2 => 
                           n8946, ZN => n9346);
   U8056 : OAI22_X1 port map( A1 => n9233, A2 => n11617, B1 => n8977, B2 => 
                           n11613, ZN => n10477);
   U8057 : OAI22_X1 port map( A1 => n9232, A2 => n11617, B1 => n8976, B2 => 
                           n11613, ZN => n10448);
   U8058 : OAI22_X1 port map( A1 => n9231, A2 => n11617, B1 => n8975, B2 => 
                           n11613, ZN => n10431);
   U8059 : OAI22_X1 port map( A1 => n9230, A2 => n11617, B1 => n8974, B2 => 
                           n11613, ZN => n10414);
   U8060 : OAI22_X1 port map( A1 => n9229, A2 => n11617, B1 => n8973, B2 => 
                           n11613, ZN => n10397);
   U8061 : OAI22_X1 port map( A1 => n9228, A2 => n11617, B1 => n8972, B2 => 
                           n11613, ZN => n10380);
   U8062 : OAI22_X1 port map( A1 => n9227, A2 => n11617, B1 => n8971, B2 => 
                           n11613, ZN => n10363);
   U8063 : OAI22_X1 port map( A1 => n9226, A2 => n11617, B1 => n8970, B2 => 
                           n11613, ZN => n10346);
   U8064 : OAI22_X1 port map( A1 => n9225, A2 => n11617, B1 => n8969, B2 => 
                           n11613, ZN => n10329);
   U8065 : OAI22_X1 port map( A1 => n9224, A2 => n11617, B1 => n8968, B2 => 
                           n11613, ZN => n10312);
   U8066 : OAI22_X1 port map( A1 => n9223, A2 => n11617, B1 => n8967, B2 => 
                           n11613, ZN => n10295);
   U8067 : OAI22_X1 port map( A1 => n9222, A2 => n11617, B1 => n8966, B2 => 
                           n11613, ZN => n10278);
   U8068 : OAI22_X1 port map( A1 => n9221, A2 => n11618, B1 => n8965, B2 => 
                           n11614, ZN => n10261);
   U8069 : OAI22_X1 port map( A1 => n9220, A2 => n11618, B1 => n8964, B2 => 
                           n11614, ZN => n10244);
   U8070 : OAI22_X1 port map( A1 => n9219, A2 => n11618, B1 => n8963, B2 => 
                           n11614, ZN => n10227);
   U8071 : OAI22_X1 port map( A1 => n9218, A2 => n11618, B1 => n8962, B2 => 
                           n11614, ZN => n10210);
   U8072 : OAI22_X1 port map( A1 => n9217, A2 => n11618, B1 => n8961, B2 => 
                           n11614, ZN => n10193);
   U8073 : OAI22_X1 port map( A1 => n9216, A2 => n11618, B1 => n8960, B2 => 
                           n11614, ZN => n10176);
   U8074 : OAI22_X1 port map( A1 => n9215, A2 => n11618, B1 => n8959, B2 => 
                           n11614, ZN => n10159);
   U8075 : OAI22_X1 port map( A1 => n9214, A2 => n11618, B1 => n8958, B2 => 
                           n11614, ZN => n10142);
   U8076 : OAI22_X1 port map( A1 => n9213, A2 => n11618, B1 => n8957, B2 => 
                           n11614, ZN => n10125);
   U8077 : OAI22_X1 port map( A1 => n9212, A2 => n11618, B1 => n8956, B2 => 
                           n11614, ZN => n10108);
   U8078 : OAI22_X1 port map( A1 => n9211, A2 => n11618, B1 => n8955, B2 => 
                           n11614, ZN => n10091);
   U8079 : OAI22_X1 port map( A1 => n9210, A2 => n11618, B1 => n8954, B2 => 
                           n11614, ZN => n10074);
   U8080 : OAI22_X1 port map( A1 => n9209, A2 => n11619, B1 => n8953, B2 => 
                           n11615, ZN => n10057);
   U8081 : OAI22_X1 port map( A1 => n9208, A2 => n11619, B1 => n8952, B2 => 
                           n11615, ZN => n10040);
   U8082 : OAI22_X1 port map( A1 => n9207, A2 => n11619, B1 => n8951, B2 => 
                           n11615, ZN => n10023);
   U8083 : OAI22_X1 port map( A1 => n9206, A2 => n11619, B1 => n8950, B2 => 
                           n11615, ZN => n10006);
   U8084 : OAI22_X1 port map( A1 => n9205, A2 => n11619, B1 => n8949, B2 => 
                           n11615, ZN => n9989);
   U8085 : OAI22_X1 port map( A1 => n9204, A2 => n11619, B1 => n8948, B2 => 
                           n11615, ZN => n9972);
   U8086 : OAI22_X1 port map( A1 => n9203, A2 => n11619, B1 => n8947, B2 => 
                           n11615, ZN => n9955);
   U8087 : OAI22_X1 port map( A1 => n9202, A2 => n11619, B1 => n8946, B2 => 
                           n11615, ZN => n9936);
   U8088 : OAI22_X1 port map( A1 => n11878, A2 => n8913, B1 => n11874, B2 => 
                           n9105, ZN => n9863);
   U8089 : OAI22_X1 port map( A1 => n11878, A2 => n8912, B1 => n11874, B2 => 
                           n9104, ZN => n9846);
   U8090 : OAI22_X1 port map( A1 => n11878, A2 => n8911, B1 => n11874, B2 => 
                           n9103, ZN => n9829);
   U8091 : OAI22_X1 port map( A1 => n11878, A2 => n8910, B1 => n11874, B2 => 
                           n9102, ZN => n9812);
   U8092 : OAI22_X1 port map( A1 => n11878, A2 => n8909, B1 => n11874, B2 => 
                           n9101, ZN => n9795);
   U8093 : OAI22_X1 port map( A1 => n11878, A2 => n8908, B1 => n11874, B2 => 
                           n9100, ZN => n9778);
   U8094 : OAI22_X1 port map( A1 => n11878, A2 => n8907, B1 => n11874, B2 => 
                           n9099, ZN => n9761);
   U8095 : OAI22_X1 port map( A1 => n11878, A2 => n8906, B1 => n11874, B2 => 
                           n9098, ZN => n9744);
   U8096 : OAI22_X1 port map( A1 => n11878, A2 => n8905, B1 => n11874, B2 => 
                           n9097, ZN => n9727);
   U8097 : OAI22_X1 port map( A1 => n11878, A2 => n8904, B1 => n11874, B2 => 
                           n9096, ZN => n9710);
   U8098 : OAI22_X1 port map( A1 => n11878, A2 => n8903, B1 => n11874, B2 => 
                           n9095, ZN => n9693);
   U8099 : OAI22_X1 port map( A1 => n11878, A2 => n8902, B1 => n11874, B2 => 
                           n9094, ZN => n9676);
   U8100 : OAI22_X1 port map( A1 => n11879, A2 => n8901, B1 => n11875, B2 => 
                           n9093, ZN => n9659);
   U8101 : OAI22_X1 port map( A1 => n11879, A2 => n8900, B1 => n11875, B2 => 
                           n9092, ZN => n9642);
   U8102 : OAI22_X1 port map( A1 => n11879, A2 => n8899, B1 => n11875, B2 => 
                           n9091, ZN => n9625);
   U8103 : OAI22_X1 port map( A1 => n11879, A2 => n8898, B1 => n11875, B2 => 
                           n9090, ZN => n9608);
   U8104 : OAI22_X1 port map( A1 => n11879, A2 => n8897, B1 => n11875, B2 => 
                           n9089, ZN => n9591);
   U8105 : OAI22_X1 port map( A1 => n11879, A2 => n8896, B1 => n11875, B2 => 
                           n9088, ZN => n9574);
   U8106 : OAI22_X1 port map( A1 => n11879, A2 => n8895, B1 => n11875, B2 => 
                           n9087, ZN => n9557);
   U8107 : OAI22_X1 port map( A1 => n11879, A2 => n8894, B1 => n11875, B2 => 
                           n9086, ZN => n9540);
   U8108 : OAI22_X1 port map( A1 => n11879, A2 => n8893, B1 => n11875, B2 => 
                           n9085, ZN => n9523);
   U8109 : OAI22_X1 port map( A1 => n11879, A2 => n8892, B1 => n11875, B2 => 
                           n9084, ZN => n9506);
   U8110 : OAI22_X1 port map( A1 => n11879, A2 => n8891, B1 => n11875, B2 => 
                           n9083, ZN => n9489);
   U8111 : OAI22_X1 port map( A1 => n11879, A2 => n8890, B1 => n11875, B2 => 
                           n9082, ZN => n9472);
   U8112 : OAI22_X1 port map( A1 => n11880, A2 => n8889, B1 => n11876, B2 => 
                           n9081, ZN => n9455);
   U8113 : OAI22_X1 port map( A1 => n11880, A2 => n8888, B1 => n11876, B2 => 
                           n9080, ZN => n9438);
   U8114 : OAI22_X1 port map( A1 => n11880, A2 => n8887, B1 => n11876, B2 => 
                           n9079, ZN => n9421);
   U8115 : OAI22_X1 port map( A1 => n11880, A2 => n8886, B1 => n11876, B2 => 
                           n9078, ZN => n9404);
   U8116 : OAI22_X1 port map( A1 => n11880, A2 => n8885, B1 => n11876, B2 => 
                           n9077, ZN => n9387);
   U8117 : OAI22_X1 port map( A1 => n11880, A2 => n8884, B1 => n11876, B2 => 
                           n9076, ZN => n9370);
   U8118 : OAI22_X1 port map( A1 => n11880, A2 => n8883, B1 => n11876, B2 => 
                           n9075, ZN => n9353);
   U8119 : OAI22_X1 port map( A1 => n11880, A2 => n8882, B1 => n11876, B2 => 
                           n9074, ZN => n9304);
   U8120 : OAI22_X1 port map( A1 => n11862, A2 => n9201, B1 => n11858, B2 => 
                           n9297, ZN => n9869);
   U8121 : OAI22_X1 port map( A1 => n11862, A2 => n9200, B1 => n11858, B2 => 
                           n9296, ZN => n9847);
   U8122 : OAI22_X1 port map( A1 => n11862, A2 => n9199, B1 => n11858, B2 => 
                           n9295, ZN => n9830);
   U8123 : OAI22_X1 port map( A1 => n11862, A2 => n9198, B1 => n11858, B2 => 
                           n9294, ZN => n9813);
   U8124 : OAI22_X1 port map( A1 => n11862, A2 => n9197, B1 => n11858, B2 => 
                           n9293, ZN => n9796);
   U8125 : OAI22_X1 port map( A1 => n11862, A2 => n9196, B1 => n11858, B2 => 
                           n9292, ZN => n9779);
   U8126 : OAI22_X1 port map( A1 => n11862, A2 => n9195, B1 => n11858, B2 => 
                           n9291, ZN => n9762);
   U8127 : OAI22_X1 port map( A1 => n11862, A2 => n9194, B1 => n11858, B2 => 
                           n9290, ZN => n9745);
   U8128 : OAI22_X1 port map( A1 => n11862, A2 => n9193, B1 => n11858, B2 => 
                           n9289, ZN => n9728);
   U8129 : OAI22_X1 port map( A1 => n11862, A2 => n9192, B1 => n11858, B2 => 
                           n9288, ZN => n9711);
   U8130 : OAI22_X1 port map( A1 => n11862, A2 => n9191, B1 => n11858, B2 => 
                           n9287, ZN => n9694);
   U8131 : OAI22_X1 port map( A1 => n11862, A2 => n9190, B1 => n11858, B2 => 
                           n9286, ZN => n9677);
   U8132 : OAI22_X1 port map( A1 => n11863, A2 => n9189, B1 => n11859, B2 => 
                           n9285, ZN => n9660);
   U8133 : OAI22_X1 port map( A1 => n11863, A2 => n9188, B1 => n11859, B2 => 
                           n9284, ZN => n9643);
   U8134 : OAI22_X1 port map( A1 => n11863, A2 => n9187, B1 => n11859, B2 => 
                           n9283, ZN => n9626);
   U8135 : OAI22_X1 port map( A1 => n11863, A2 => n9186, B1 => n11859, B2 => 
                           n9282, ZN => n9609);
   U8136 : OAI22_X1 port map( A1 => n11863, A2 => n9185, B1 => n11859, B2 => 
                           n9281, ZN => n9592);
   U8137 : OAI22_X1 port map( A1 => n11863, A2 => n9184, B1 => n11859, B2 => 
                           n9280, ZN => n9575);
   U8138 : OAI22_X1 port map( A1 => n11863, A2 => n9183, B1 => n11859, B2 => 
                           n9279, ZN => n9558);
   U8139 : OAI22_X1 port map( A1 => n11863, A2 => n9182, B1 => n11859, B2 => 
                           n9278, ZN => n9541);
   U8140 : OAI22_X1 port map( A1 => n11863, A2 => n9181, B1 => n11859, B2 => 
                           n9277, ZN => n9524);
   U8141 : OAI22_X1 port map( A1 => n11863, A2 => n9180, B1 => n11859, B2 => 
                           n9276, ZN => n9507);
   U8142 : OAI22_X1 port map( A1 => n11863, A2 => n9179, B1 => n11859, B2 => 
                           n9275, ZN => n9490);
   U8143 : OAI22_X1 port map( A1 => n11863, A2 => n9178, B1 => n11859, B2 => 
                           n9274, ZN => n9473);
   U8144 : OAI22_X1 port map( A1 => n11864, A2 => n9177, B1 => n11860, B2 => 
                           n9273, ZN => n9456);
   U8145 : OAI22_X1 port map( A1 => n11864, A2 => n9176, B1 => n11860, B2 => 
                           n9272, ZN => n9439);
   U8146 : OAI22_X1 port map( A1 => n11864, A2 => n9175, B1 => n11860, B2 => 
                           n9271, ZN => n9422);
   U8147 : OAI22_X1 port map( A1 => n11864, A2 => n9174, B1 => n11860, B2 => 
                           n9270, ZN => n9405);
   U8148 : OAI22_X1 port map( A1 => n11864, A2 => n9173, B1 => n11860, B2 => 
                           n9269, ZN => n9388);
   U8149 : OAI22_X1 port map( A1 => n11864, A2 => n9172, B1 => n11860, B2 => 
                           n9268, ZN => n9371);
   U8150 : OAI22_X1 port map( A1 => n11864, A2 => n9171, B1 => n11860, B2 => 
                           n9267, ZN => n9354);
   U8151 : OAI22_X1 port map( A1 => n11864, A2 => n9170, B1 => n11860, B2 => 
                           n9266, ZN => n9309);
   U8152 : OAI22_X1 port map( A1 => n8913, A2 => n11739, B1 => n9105, B2 => 
                           n11735, ZN => n10453);
   U8153 : OAI22_X1 port map( A1 => n8912, A2 => n11739, B1 => n9104, B2 => 
                           n11735, ZN => n10436);
   U8154 : OAI22_X1 port map( A1 => n8911, A2 => n11739, B1 => n9103, B2 => 
                           n11735, ZN => n10419);
   U8155 : OAI22_X1 port map( A1 => n8910, A2 => n11739, B1 => n9102, B2 => 
                           n11735, ZN => n10402);
   U8156 : OAI22_X1 port map( A1 => n8909, A2 => n11739, B1 => n9101, B2 => 
                           n11735, ZN => n10385);
   U8157 : OAI22_X1 port map( A1 => n8908, A2 => n11739, B1 => n9100, B2 => 
                           n11735, ZN => n10368);
   U8158 : OAI22_X1 port map( A1 => n8907, A2 => n11739, B1 => n9099, B2 => 
                           n11735, ZN => n10351);
   U8159 : OAI22_X1 port map( A1 => n8906, A2 => n11739, B1 => n9098, B2 => 
                           n11735, ZN => n10334);
   U8160 : OAI22_X1 port map( A1 => n8905, A2 => n11739, B1 => n9097, B2 => 
                           n11735, ZN => n10317);
   U8161 : OAI22_X1 port map( A1 => n8904, A2 => n11739, B1 => n9096, B2 => 
                           n11735, ZN => n10300);
   U8162 : OAI22_X1 port map( A1 => n8903, A2 => n11739, B1 => n9095, B2 => 
                           n11735, ZN => n10283);
   U8163 : OAI22_X1 port map( A1 => n8902, A2 => n11739, B1 => n9094, B2 => 
                           n11735, ZN => n10266);
   U8164 : OAI22_X1 port map( A1 => n8901, A2 => n11740, B1 => n9093, B2 => 
                           n11736, ZN => n10249);
   U8165 : OAI22_X1 port map( A1 => n8900, A2 => n11740, B1 => n9092, B2 => 
                           n11736, ZN => n10232);
   U8166 : OAI22_X1 port map( A1 => n8899, A2 => n11740, B1 => n9091, B2 => 
                           n11736, ZN => n10215);
   U8167 : OAI22_X1 port map( A1 => n8898, A2 => n11740, B1 => n9090, B2 => 
                           n11736, ZN => n10198);
   U8168 : OAI22_X1 port map( A1 => n8897, A2 => n11740, B1 => n9089, B2 => 
                           n11736, ZN => n10181);
   U8169 : OAI22_X1 port map( A1 => n8896, A2 => n11740, B1 => n9088, B2 => 
                           n11736, ZN => n10164);
   U8170 : OAI22_X1 port map( A1 => n8895, A2 => n11740, B1 => n9087, B2 => 
                           n11736, ZN => n10147);
   U8171 : OAI22_X1 port map( A1 => n8894, A2 => n11740, B1 => n9086, B2 => 
                           n11736, ZN => n10130);
   U8172 : OAI22_X1 port map( A1 => n8893, A2 => n11740, B1 => n9085, B2 => 
                           n11736, ZN => n10113);
   U8173 : OAI22_X1 port map( A1 => n8892, A2 => n11740, B1 => n9084, B2 => 
                           n11736, ZN => n10096);
   U8174 : OAI22_X1 port map( A1 => n8891, A2 => n11740, B1 => n9083, B2 => 
                           n11736, ZN => n10079);
   U8175 : OAI22_X1 port map( A1 => n8890, A2 => n11740, B1 => n9082, B2 => 
                           n11736, ZN => n10062);
   U8176 : OAI22_X1 port map( A1 => n8889, A2 => n11741, B1 => n9081, B2 => 
                           n11737, ZN => n10045);
   U8177 : OAI22_X1 port map( A1 => n8888, A2 => n11741, B1 => n9080, B2 => 
                           n11737, ZN => n10028);
   U8178 : OAI22_X1 port map( A1 => n8887, A2 => n11741, B1 => n9079, B2 => 
                           n11737, ZN => n10011);
   U8179 : OAI22_X1 port map( A1 => n8886, A2 => n11741, B1 => n9078, B2 => 
                           n11737, ZN => n9994);
   U8180 : OAI22_X1 port map( A1 => n8885, A2 => n11741, B1 => n9077, B2 => 
                           n11737, ZN => n9977);
   U8181 : OAI22_X1 port map( A1 => n8884, A2 => n11741, B1 => n9076, B2 => 
                           n11737, ZN => n9960);
   U8182 : OAI22_X1 port map( A1 => n8883, A2 => n11741, B1 => n9075, B2 => 
                           n11737, ZN => n9943);
   U8183 : OAI22_X1 port map( A1 => n8882, A2 => n11741, B1 => n9074, B2 => 
                           n11737, ZN => n9894);
   U8184 : OAI22_X1 port map( A1 => n11846, A2 => n8881, B1 => n11842, B2 => 
                           n8945, ZN => n9872);
   U8185 : OAI22_X1 port map( A1 => n11846, A2 => n8880, B1 => n11842, B2 => 
                           n8944, ZN => n9848);
   U8186 : OAI22_X1 port map( A1 => n11846, A2 => n8879, B1 => n11842, B2 => 
                           n8943, ZN => n9831);
   U8187 : OAI22_X1 port map( A1 => n11846, A2 => n8878, B1 => n11842, B2 => 
                           n8942, ZN => n9814);
   U8188 : OAI22_X1 port map( A1 => n11846, A2 => n8877, B1 => n11842, B2 => 
                           n8941, ZN => n9797);
   U8189 : OAI22_X1 port map( A1 => n11846, A2 => n8876, B1 => n11842, B2 => 
                           n8940, ZN => n9780);
   U8190 : OAI22_X1 port map( A1 => n11846, A2 => n8875, B1 => n11842, B2 => 
                           n8939, ZN => n9763);
   U8191 : OAI22_X1 port map( A1 => n11846, A2 => n8874, B1 => n11842, B2 => 
                           n8938, ZN => n9746);
   U8192 : OAI22_X1 port map( A1 => n11846, A2 => n8873, B1 => n11842, B2 => 
                           n8937, ZN => n9729);
   U8193 : OAI22_X1 port map( A1 => n11846, A2 => n8872, B1 => n11842, B2 => 
                           n8936, ZN => n9712);
   U8194 : OAI22_X1 port map( A1 => n11846, A2 => n8871, B1 => n11842, B2 => 
                           n8935, ZN => n9695);
   U8195 : OAI22_X1 port map( A1 => n11846, A2 => n8870, B1 => n11842, B2 => 
                           n8934, ZN => n9678);
   U8196 : OAI22_X1 port map( A1 => n11847, A2 => n8869, B1 => n11843, B2 => 
                           n8933, ZN => n9661);
   U8197 : OAI22_X1 port map( A1 => n11847, A2 => n8868, B1 => n11843, B2 => 
                           n8932, ZN => n9644);
   U8198 : OAI22_X1 port map( A1 => n11847, A2 => n8867, B1 => n11843, B2 => 
                           n8931, ZN => n9627);
   U8199 : OAI22_X1 port map( A1 => n11847, A2 => n8866, B1 => n11843, B2 => 
                           n8930, ZN => n9610);
   U8200 : OAI22_X1 port map( A1 => n11847, A2 => n8865, B1 => n11843, B2 => 
                           n8929, ZN => n9593);
   U8201 : OAI22_X1 port map( A1 => n11847, A2 => n8864, B1 => n11843, B2 => 
                           n8928, ZN => n9576);
   U8202 : OAI22_X1 port map( A1 => n11847, A2 => n8863, B1 => n11843, B2 => 
                           n8927, ZN => n9559);
   U8203 : OAI22_X1 port map( A1 => n11847, A2 => n8862, B1 => n11843, B2 => 
                           n8926, ZN => n9542);
   U8204 : OAI22_X1 port map( A1 => n11847, A2 => n8861, B1 => n11843, B2 => 
                           n8925, ZN => n9525);
   U8205 : OAI22_X1 port map( A1 => n11847, A2 => n8860, B1 => n11843, B2 => 
                           n8924, ZN => n9508);
   U8206 : OAI22_X1 port map( A1 => n11847, A2 => n8859, B1 => n11843, B2 => 
                           n8923, ZN => n9491);
   U8207 : OAI22_X1 port map( A1 => n11847, A2 => n8858, B1 => n11843, B2 => 
                           n8922, ZN => n9474);
   U8208 : OAI22_X1 port map( A1 => n11848, A2 => n8857, B1 => n11844, B2 => 
                           n8921, ZN => n9457);
   U8209 : OAI22_X1 port map( A1 => n11848, A2 => n8856, B1 => n11844, B2 => 
                           n8920, ZN => n9440);
   U8210 : OAI22_X1 port map( A1 => n11848, A2 => n8855, B1 => n11844, B2 => 
                           n8919, ZN => n9423);
   U8211 : OAI22_X1 port map( A1 => n11848, A2 => n8854, B1 => n11844, B2 => 
                           n8918, ZN => n9406);
   U8212 : OAI22_X1 port map( A1 => n11848, A2 => n8853, B1 => n11844, B2 => 
                           n8917, ZN => n9389);
   U8213 : OAI22_X1 port map( A1 => n11848, A2 => n8852, B1 => n11844, B2 => 
                           n8916, ZN => n9372);
   U8214 : OAI22_X1 port map( A1 => n11848, A2 => n8851, B1 => n11844, B2 => 
                           n8915, ZN => n9355);
   U8215 : OAI22_X1 port map( A1 => n11848, A2 => n8850, B1 => n11844, B2 => 
                           n8914, ZN => n9314);
   U8216 : OAI22_X1 port map( A1 => n9201, A2 => n11723, B1 => n9297, B2 => 
                           n11719, ZN => n10459);
   U8217 : OAI22_X1 port map( A1 => n9200, A2 => n11723, B1 => n9296, B2 => 
                           n11719, ZN => n10437);
   U8218 : OAI22_X1 port map( A1 => n9199, A2 => n11723, B1 => n9295, B2 => 
                           n11719, ZN => n10420);
   U8219 : OAI22_X1 port map( A1 => n9198, A2 => n11723, B1 => n9294, B2 => 
                           n11719, ZN => n10403);
   U8220 : OAI22_X1 port map( A1 => n9197, A2 => n11723, B1 => n9293, B2 => 
                           n11719, ZN => n10386);
   U8221 : OAI22_X1 port map( A1 => n9196, A2 => n11723, B1 => n9292, B2 => 
                           n11719, ZN => n10369);
   U8222 : OAI22_X1 port map( A1 => n9195, A2 => n11723, B1 => n9291, B2 => 
                           n11719, ZN => n10352);
   U8223 : OAI22_X1 port map( A1 => n9194, A2 => n11723, B1 => n9290, B2 => 
                           n11719, ZN => n10335);
   U8224 : OAI22_X1 port map( A1 => n9193, A2 => n11723, B1 => n9289, B2 => 
                           n11719, ZN => n10318);
   U8225 : OAI22_X1 port map( A1 => n9192, A2 => n11723, B1 => n9288, B2 => 
                           n11719, ZN => n10301);
   U8226 : OAI22_X1 port map( A1 => n9191, A2 => n11723, B1 => n9287, B2 => 
                           n11719, ZN => n10284);
   U8227 : OAI22_X1 port map( A1 => n9190, A2 => n11723, B1 => n9286, B2 => 
                           n11719, ZN => n10267);
   U8228 : OAI22_X1 port map( A1 => n9189, A2 => n11724, B1 => n9285, B2 => 
                           n11720, ZN => n10250);
   U8229 : OAI22_X1 port map( A1 => n9188, A2 => n11724, B1 => n9284, B2 => 
                           n11720, ZN => n10233);
   U8230 : OAI22_X1 port map( A1 => n9187, A2 => n11724, B1 => n9283, B2 => 
                           n11720, ZN => n10216);
   U8231 : OAI22_X1 port map( A1 => n9186, A2 => n11724, B1 => n9282, B2 => 
                           n11720, ZN => n10199);
   U8232 : OAI22_X1 port map( A1 => n9185, A2 => n11724, B1 => n9281, B2 => 
                           n11720, ZN => n10182);
   U8233 : OAI22_X1 port map( A1 => n9184, A2 => n11724, B1 => n9280, B2 => 
                           n11720, ZN => n10165);
   U8234 : OAI22_X1 port map( A1 => n9183, A2 => n11724, B1 => n9279, B2 => 
                           n11720, ZN => n10148);
   U8235 : OAI22_X1 port map( A1 => n9182, A2 => n11724, B1 => n9278, B2 => 
                           n11720, ZN => n10131);
   U8236 : OAI22_X1 port map( A1 => n9181, A2 => n11724, B1 => n9277, B2 => 
                           n11720, ZN => n10114);
   U8237 : OAI22_X1 port map( A1 => n9180, A2 => n11724, B1 => n9276, B2 => 
                           n11720, ZN => n10097);
   U8238 : OAI22_X1 port map( A1 => n9179, A2 => n11724, B1 => n9275, B2 => 
                           n11720, ZN => n10080);
   U8239 : OAI22_X1 port map( A1 => n9178, A2 => n11724, B1 => n9274, B2 => 
                           n11720, ZN => n10063);
   U8240 : OAI22_X1 port map( A1 => n9177, A2 => n11725, B1 => n9273, B2 => 
                           n11721, ZN => n10046);
   U8241 : OAI22_X1 port map( A1 => n9176, A2 => n11725, B1 => n9272, B2 => 
                           n11721, ZN => n10029);
   U8242 : OAI22_X1 port map( A1 => n9175, A2 => n11725, B1 => n9271, B2 => 
                           n11721, ZN => n10012);
   U8243 : OAI22_X1 port map( A1 => n9174, A2 => n11725, B1 => n9270, B2 => 
                           n11721, ZN => n9995);
   U8244 : OAI22_X1 port map( A1 => n9173, A2 => n11725, B1 => n9269, B2 => 
                           n11721, ZN => n9978);
   U8245 : OAI22_X1 port map( A1 => n9172, A2 => n11725, B1 => n9268, B2 => 
                           n11721, ZN => n9961);
   U8246 : OAI22_X1 port map( A1 => n9171, A2 => n11725, B1 => n9267, B2 => 
                           n11721, ZN => n9944);
   U8247 : OAI22_X1 port map( A1 => n9170, A2 => n11725, B1 => n9266, B2 => 
                           n11721, ZN => n9899);
   U8248 : OAI22_X1 port map( A1 => n8881, A2 => n11707, B1 => n8945, B2 => 
                           n11703, ZN => n10462);
   U8249 : OAI22_X1 port map( A1 => n8880, A2 => n11707, B1 => n8944, B2 => 
                           n11703, ZN => n10438);
   U8250 : OAI22_X1 port map( A1 => n8879, A2 => n11707, B1 => n8943, B2 => 
                           n11703, ZN => n10421);
   U8251 : OAI22_X1 port map( A1 => n8878, A2 => n11707, B1 => n8942, B2 => 
                           n11703, ZN => n10404);
   U8252 : OAI22_X1 port map( A1 => n8877, A2 => n11707, B1 => n8941, B2 => 
                           n11703, ZN => n10387);
   U8253 : OAI22_X1 port map( A1 => n8876, A2 => n11707, B1 => n8940, B2 => 
                           n11703, ZN => n10370);
   U8254 : OAI22_X1 port map( A1 => n8875, A2 => n11707, B1 => n8939, B2 => 
                           n11703, ZN => n10353);
   U8255 : OAI22_X1 port map( A1 => n8874, A2 => n11707, B1 => n8938, B2 => 
                           n11703, ZN => n10336);
   U8256 : OAI22_X1 port map( A1 => n8873, A2 => n11707, B1 => n8937, B2 => 
                           n11703, ZN => n10319);
   U8257 : OAI22_X1 port map( A1 => n8872, A2 => n11707, B1 => n8936, B2 => 
                           n11703, ZN => n10302);
   U8258 : OAI22_X1 port map( A1 => n8871, A2 => n11707, B1 => n8935, B2 => 
                           n11703, ZN => n10285);
   U8259 : OAI22_X1 port map( A1 => n8870, A2 => n11707, B1 => n8934, B2 => 
                           n11703, ZN => n10268);
   U8260 : OAI22_X1 port map( A1 => n8869, A2 => n11708, B1 => n8933, B2 => 
                           n11704, ZN => n10251);
   U8261 : OAI22_X1 port map( A1 => n8868, A2 => n11708, B1 => n8932, B2 => 
                           n11704, ZN => n10234);
   U8262 : OAI22_X1 port map( A1 => n8867, A2 => n11708, B1 => n8931, B2 => 
                           n11704, ZN => n10217);
   U8263 : OAI22_X1 port map( A1 => n8866, A2 => n11708, B1 => n8930, B2 => 
                           n11704, ZN => n10200);
   U8264 : OAI22_X1 port map( A1 => n8865, A2 => n11708, B1 => n8929, B2 => 
                           n11704, ZN => n10183);
   U8265 : OAI22_X1 port map( A1 => n8864, A2 => n11708, B1 => n8928, B2 => 
                           n11704, ZN => n10166);
   U8266 : OAI22_X1 port map( A1 => n8863, A2 => n11708, B1 => n8927, B2 => 
                           n11704, ZN => n10149);
   U8267 : OAI22_X1 port map( A1 => n8862, A2 => n11708, B1 => n8926, B2 => 
                           n11704, ZN => n10132);
   U8268 : OAI22_X1 port map( A1 => n8861, A2 => n11708, B1 => n8925, B2 => 
                           n11704, ZN => n10115);
   U8269 : OAI22_X1 port map( A1 => n8860, A2 => n11708, B1 => n8924, B2 => 
                           n11704, ZN => n10098);
   U8270 : OAI22_X1 port map( A1 => n8859, A2 => n11708, B1 => n8923, B2 => 
                           n11704, ZN => n10081);
   U8271 : OAI22_X1 port map( A1 => n8858, A2 => n11708, B1 => n8922, B2 => 
                           n11704, ZN => n10064);
   U8272 : OAI22_X1 port map( A1 => n8857, A2 => n11709, B1 => n8921, B2 => 
                           n11705, ZN => n10047);
   U8273 : OAI22_X1 port map( A1 => n8856, A2 => n11709, B1 => n8920, B2 => 
                           n11705, ZN => n10030);
   U8274 : OAI22_X1 port map( A1 => n8855, A2 => n11709, B1 => n8919, B2 => 
                           n11705, ZN => n10013);
   U8275 : OAI22_X1 port map( A1 => n8854, A2 => n11709, B1 => n8918, B2 => 
                           n11705, ZN => n9996);
   U8276 : OAI22_X1 port map( A1 => n8853, A2 => n11709, B1 => n8917, B2 => 
                           n11705, ZN => n9979);
   U8277 : OAI22_X1 port map( A1 => n8852, A2 => n11709, B1 => n8916, B2 => 
                           n11705, ZN => n9962);
   U8278 : OAI22_X1 port map( A1 => n8851, A2 => n11709, B1 => n8915, B2 => 
                           n11705, ZN => n9945);
   U8279 : OAI22_X1 port map( A1 => n8850, A2 => n11709, B1 => n8914, B2 => 
                           n11705, ZN => n9904);
   U8280 : OAI22_X1 port map( A1 => n11268, A2 => n11483, B1 => n9233, B2 => 
                           n11364, ZN => n1342);
   U8281 : OAI22_X1 port map( A1 => n11268, A2 => n11487, B1 => n9232, B2 => 
                           n11364, ZN => n1343);
   U8282 : OAI22_X1 port map( A1 => n11268, A2 => n11491, B1 => n9231, B2 => 
                           n11364, ZN => n1344);
   U8283 : OAI22_X1 port map( A1 => n11268, A2 => n11495, B1 => n9230, B2 => 
                           n11364, ZN => n1345);
   U8284 : OAI22_X1 port map( A1 => n11268, A2 => n11499, B1 => n9229, B2 => 
                           n11364, ZN => n1346);
   U8285 : OAI22_X1 port map( A1 => n11268, A2 => n11503, B1 => n9228, B2 => 
                           n11364, ZN => n1347);
   U8286 : OAI22_X1 port map( A1 => n11268, A2 => n11507, B1 => n9227, B2 => 
                           n11364, ZN => n1348);
   U8287 : OAI22_X1 port map( A1 => n11268, A2 => n11511, B1 => n9226, B2 => 
                           n11364, ZN => n1349);
   U8288 : OAI22_X1 port map( A1 => n11267, A2 => n11515, B1 => n9225, B2 => 
                           n11364, ZN => n1350);
   U8289 : OAI22_X1 port map( A1 => n11267, A2 => n11519, B1 => n9224, B2 => 
                           n11364, ZN => n1351);
   U8290 : OAI22_X1 port map( A1 => n11267, A2 => n11523, B1 => n9223, B2 => 
                           n11364, ZN => n1352);
   U8291 : OAI22_X1 port map( A1 => n11267, A2 => n11527, B1 => n9222, B2 => 
                           n11364, ZN => n1353);
   U8292 : OAI22_X1 port map( A1 => n11267, A2 => n11531, B1 => n9221, B2 => 
                           n10553, ZN => n1354);
   U8293 : OAI22_X1 port map( A1 => n11267, A2 => n11535, B1 => n9220, B2 => 
                           n10553, ZN => n1355);
   U8294 : OAI22_X1 port map( A1 => n11267, A2 => n11539, B1 => n9219, B2 => 
                           n10553, ZN => n1356);
   U8295 : OAI22_X1 port map( A1 => n11267, A2 => n11543, B1 => n9218, B2 => 
                           n11364, ZN => n1357);
   U8296 : OAI22_X1 port map( A1 => n11267, A2 => n11547, B1 => n9217, B2 => 
                           n11364, ZN => n1358);
   U8297 : OAI22_X1 port map( A1 => n11267, A2 => n11551, B1 => n9216, B2 => 
                           n11364, ZN => n1359);
   U8298 : OAI22_X1 port map( A1 => n11267, A2 => n11555, B1 => n9215, B2 => 
                           n11364, ZN => n1360);
   U8299 : OAI22_X1 port map( A1 => n11267, A2 => n11559, B1 => n9214, B2 => 
                           n11364, ZN => n1361);
   U8300 : OAI22_X1 port map( A1 => n11266, A2 => n11563, B1 => n9213, B2 => 
                           n11364, ZN => n1362);
   U8301 : OAI22_X1 port map( A1 => n11266, A2 => n11567, B1 => n9212, B2 => 
                           n11364, ZN => n1363);
   U8302 : OAI22_X1 port map( A1 => n11266, A2 => n11571, B1 => n9211, B2 => 
                           n11364, ZN => n1364);
   U8303 : OAI22_X1 port map( A1 => n11266, A2 => n11575, B1 => n9210, B2 => 
                           n11364, ZN => n1365);
   U8304 : OAI22_X1 port map( A1 => n11266, A2 => n11579, B1 => n9209, B2 => 
                           n10553, ZN => n1366);
   U8305 : OAI22_X1 port map( A1 => n11266, A2 => n11583, B1 => n9208, B2 => 
                           n10553, ZN => n1367);
   U8306 : OAI22_X1 port map( A1 => n11266, A2 => n11587, B1 => n9207, B2 => 
                           n10553, ZN => n1368);
   U8307 : OAI22_X1 port map( A1 => n11266, A2 => n11591, B1 => n9206, B2 => 
                           n10553, ZN => n1369);
   U8308 : OAI22_X1 port map( A1 => n11266, A2 => n11595, B1 => n9205, B2 => 
                           n10553, ZN => n1370);
   U8309 : OAI22_X1 port map( A1 => n11266, A2 => n11599, B1 => n9204, B2 => 
                           n10553, ZN => n1371);
   U8310 : OAI22_X1 port map( A1 => n11266, A2 => n11603, B1 => n9203, B2 => 
                           n10553, ZN => n1372);
   U8311 : OAI22_X1 port map( A1 => n11266, A2 => n11611, B1 => n9202, B2 => 
                           n10553, ZN => n1373);
   U8312 : OAI22_X1 port map( A1 => n11271, A2 => n11483, B1 => n9201, B2 => 
                           n11368, ZN => n1374);
   U8313 : OAI22_X1 port map( A1 => n11271, A2 => n11487, B1 => n9200, B2 => 
                           n11368, ZN => n1375);
   U8314 : OAI22_X1 port map( A1 => n11271, A2 => n11491, B1 => n9199, B2 => 
                           n11368, ZN => n1376);
   U8315 : OAI22_X1 port map( A1 => n11271, A2 => n11495, B1 => n9198, B2 => 
                           n11368, ZN => n1377);
   U8316 : OAI22_X1 port map( A1 => n11271, A2 => n11499, B1 => n9197, B2 => 
                           n11368, ZN => n1378);
   U8317 : OAI22_X1 port map( A1 => n11271, A2 => n11503, B1 => n9196, B2 => 
                           n11368, ZN => n1379);
   U8318 : OAI22_X1 port map( A1 => n11271, A2 => n11507, B1 => n9195, B2 => 
                           n11368, ZN => n1380);
   U8319 : OAI22_X1 port map( A1 => n11271, A2 => n11511, B1 => n9194, B2 => 
                           n11368, ZN => n1381);
   U8320 : OAI22_X1 port map( A1 => n11270, A2 => n11515, B1 => n9193, B2 => 
                           n11368, ZN => n1382);
   U8321 : OAI22_X1 port map( A1 => n11270, A2 => n11519, B1 => n9192, B2 => 
                           n11368, ZN => n1383);
   U8322 : OAI22_X1 port map( A1 => n11270, A2 => n11523, B1 => n9191, B2 => 
                           n11368, ZN => n1384);
   U8323 : OAI22_X1 port map( A1 => n11270, A2 => n11527, B1 => n9190, B2 => 
                           n11368, ZN => n1385);
   U8324 : OAI22_X1 port map( A1 => n11270, A2 => n11531, B1 => n9189, B2 => 
                           n10551, ZN => n1386);
   U8325 : OAI22_X1 port map( A1 => n11270, A2 => n11535, B1 => n9188, B2 => 
                           n10551, ZN => n1387);
   U8326 : OAI22_X1 port map( A1 => n11270, A2 => n11539, B1 => n9187, B2 => 
                           n10551, ZN => n1388);
   U8327 : OAI22_X1 port map( A1 => n11270, A2 => n11543, B1 => n9186, B2 => 
                           n11368, ZN => n1389);
   U8328 : OAI22_X1 port map( A1 => n11270, A2 => n11547, B1 => n9185, B2 => 
                           n11368, ZN => n1390);
   U8329 : OAI22_X1 port map( A1 => n11270, A2 => n11551, B1 => n9184, B2 => 
                           n11368, ZN => n1391);
   U8330 : OAI22_X1 port map( A1 => n11270, A2 => n11555, B1 => n9183, B2 => 
                           n11368, ZN => n1392);
   U8331 : OAI22_X1 port map( A1 => n11270, A2 => n11559, B1 => n9182, B2 => 
                           n11368, ZN => n1393);
   U8332 : OAI22_X1 port map( A1 => n11269, A2 => n11563, B1 => n9181, B2 => 
                           n11368, ZN => n1394);
   U8333 : OAI22_X1 port map( A1 => n11269, A2 => n11567, B1 => n9180, B2 => 
                           n11368, ZN => n1395);
   U8334 : OAI22_X1 port map( A1 => n11269, A2 => n11571, B1 => n9179, B2 => 
                           n11368, ZN => n1396);
   U8335 : OAI22_X1 port map( A1 => n11269, A2 => n11575, B1 => n9178, B2 => 
                           n11368, ZN => n1397);
   U8336 : OAI22_X1 port map( A1 => n11269, A2 => n11579, B1 => n9177, B2 => 
                           n10551, ZN => n1398);
   U8337 : OAI22_X1 port map( A1 => n11269, A2 => n11583, B1 => n9176, B2 => 
                           n10551, ZN => n1399);
   U8338 : OAI22_X1 port map( A1 => n11269, A2 => n11587, B1 => n9175, B2 => 
                           n10551, ZN => n1400);
   U8339 : OAI22_X1 port map( A1 => n11269, A2 => n11591, B1 => n9174, B2 => 
                           n10551, ZN => n1401);
   U8340 : OAI22_X1 port map( A1 => n11269, A2 => n11595, B1 => n9173, B2 => 
                           n10551, ZN => n1402);
   U8341 : OAI22_X1 port map( A1 => n11269, A2 => n11599, B1 => n9172, B2 => 
                           n10551, ZN => n1403);
   U8342 : OAI22_X1 port map( A1 => n11269, A2 => n11603, B1 => n9171, B2 => 
                           n10551, ZN => n1404);
   U8343 : OAI22_X1 port map( A1 => n11269, A2 => n11611, B1 => n9170, B2 => 
                           n10551, ZN => n1405);
   U8344 : OAI22_X1 port map( A1 => n11298, A2 => n11482, B1 => n8913, B2 => 
                           n11404, ZN => n1662);
   U8345 : OAI22_X1 port map( A1 => n11298, A2 => n11486, B1 => n8912, B2 => 
                           n11404, ZN => n1663);
   U8346 : OAI22_X1 port map( A1 => n11298, A2 => n11490, B1 => n8911, B2 => 
                           n11404, ZN => n1664);
   U8347 : OAI22_X1 port map( A1 => n11298, A2 => n11494, B1 => n8910, B2 => 
                           n11404, ZN => n1665);
   U8348 : OAI22_X1 port map( A1 => n11298, A2 => n11498, B1 => n8909, B2 => 
                           n11404, ZN => n1666);
   U8349 : OAI22_X1 port map( A1 => n11298, A2 => n11502, B1 => n8908, B2 => 
                           n11404, ZN => n1667);
   U8350 : OAI22_X1 port map( A1 => n11298, A2 => n11506, B1 => n8907, B2 => 
                           n11404, ZN => n1668);
   U8351 : OAI22_X1 port map( A1 => n11298, A2 => n11510, B1 => n8906, B2 => 
                           n11404, ZN => n1669);
   U8352 : OAI22_X1 port map( A1 => n11297, A2 => n11514, B1 => n8905, B2 => 
                           n11404, ZN => n1670);
   U8353 : OAI22_X1 port map( A1 => n11297, A2 => n11518, B1 => n8904, B2 => 
                           n11404, ZN => n1671);
   U8354 : OAI22_X1 port map( A1 => n11297, A2 => n11522, B1 => n8903, B2 => 
                           n11404, ZN => n1672);
   U8355 : OAI22_X1 port map( A1 => n11297, A2 => n11526, B1 => n8902, B2 => 
                           n11404, ZN => n1673);
   U8356 : OAI22_X1 port map( A1 => n11297, A2 => n11530, B1 => n8901, B2 => 
                           n10539, ZN => n1674);
   U8357 : OAI22_X1 port map( A1 => n11297, A2 => n11534, B1 => n8900, B2 => 
                           n10539, ZN => n1675);
   U8358 : OAI22_X1 port map( A1 => n11297, A2 => n11538, B1 => n8899, B2 => 
                           n10539, ZN => n1676);
   U8359 : OAI22_X1 port map( A1 => n11297, A2 => n11542, B1 => n8898, B2 => 
                           n11404, ZN => n1677);
   U8360 : OAI22_X1 port map( A1 => n11297, A2 => n11546, B1 => n8897, B2 => 
                           n11404, ZN => n1678);
   U8361 : OAI22_X1 port map( A1 => n11297, A2 => n11550, B1 => n8896, B2 => 
                           n11404, ZN => n1679);
   U8362 : OAI22_X1 port map( A1 => n11297, A2 => n11554, B1 => n8895, B2 => 
                           n11404, ZN => n1680);
   U8363 : OAI22_X1 port map( A1 => n11297, A2 => n11558, B1 => n8894, B2 => 
                           n11404, ZN => n1681);
   U8364 : OAI22_X1 port map( A1 => n11296, A2 => n11562, B1 => n8893, B2 => 
                           n11404, ZN => n1682);
   U8365 : OAI22_X1 port map( A1 => n11296, A2 => n11566, B1 => n8892, B2 => 
                           n11404, ZN => n1683);
   U8366 : OAI22_X1 port map( A1 => n11296, A2 => n11570, B1 => n8891, B2 => 
                           n11404, ZN => n1684);
   U8367 : OAI22_X1 port map( A1 => n11296, A2 => n11574, B1 => n8890, B2 => 
                           n11404, ZN => n1685);
   U8368 : OAI22_X1 port map( A1 => n11296, A2 => n11578, B1 => n8889, B2 => 
                           n10539, ZN => n1686);
   U8369 : OAI22_X1 port map( A1 => n11296, A2 => n11582, B1 => n8888, B2 => 
                           n10539, ZN => n1687);
   U8370 : OAI22_X1 port map( A1 => n11296, A2 => n11586, B1 => n8887, B2 => 
                           n10539, ZN => n1688);
   U8371 : OAI22_X1 port map( A1 => n11296, A2 => n11590, B1 => n8886, B2 => 
                           n10539, ZN => n1689);
   U8372 : OAI22_X1 port map( A1 => n11296, A2 => n11594, B1 => n8885, B2 => 
                           n10539, ZN => n1690);
   U8373 : OAI22_X1 port map( A1 => n11296, A2 => n11598, B1 => n8884, B2 => 
                           n10539, ZN => n1691);
   U8374 : OAI22_X1 port map( A1 => n11296, A2 => n11602, B1 => n8883, B2 => 
                           n10539, ZN => n1692);
   U8375 : OAI22_X1 port map( A1 => n11296, A2 => n11610, B1 => n8882, B2 => 
                           n10539, ZN => n1693);
   U8376 : OAI22_X1 port map( A1 => n11301, A2 => n11482, B1 => n8881, B2 => 
                           n11408, ZN => n1694);
   U8377 : OAI22_X1 port map( A1 => n11301, A2 => n11486, B1 => n8880, B2 => 
                           n11408, ZN => n1695);
   U8378 : OAI22_X1 port map( A1 => n11301, A2 => n11490, B1 => n8879, B2 => 
                           n11408, ZN => n1696);
   U8379 : OAI22_X1 port map( A1 => n11301, A2 => n11494, B1 => n8878, B2 => 
                           n11408, ZN => n1697);
   U8380 : OAI22_X1 port map( A1 => n11301, A2 => n11498, B1 => n8877, B2 => 
                           n11408, ZN => n1698);
   U8381 : OAI22_X1 port map( A1 => n11301, A2 => n11502, B1 => n8876, B2 => 
                           n11408, ZN => n1699);
   U8382 : OAI22_X1 port map( A1 => n11301, A2 => n11506, B1 => n8875, B2 => 
                           n11408, ZN => n1700);
   U8383 : OAI22_X1 port map( A1 => n11301, A2 => n11510, B1 => n8874, B2 => 
                           n11408, ZN => n1701);
   U8384 : OAI22_X1 port map( A1 => n11300, A2 => n11514, B1 => n8873, B2 => 
                           n11408, ZN => n1702);
   U8385 : OAI22_X1 port map( A1 => n11300, A2 => n11518, B1 => n8872, B2 => 
                           n11408, ZN => n1703);
   U8386 : OAI22_X1 port map( A1 => n11300, A2 => n11522, B1 => n8871, B2 => 
                           n11408, ZN => n1704);
   U8387 : OAI22_X1 port map( A1 => n11300, A2 => n11526, B1 => n8870, B2 => 
                           n11408, ZN => n1705);
   U8388 : OAI22_X1 port map( A1 => n11300, A2 => n11530, B1 => n8869, B2 => 
                           n10538, ZN => n1706);
   U8389 : OAI22_X1 port map( A1 => n11300, A2 => n11534, B1 => n8868, B2 => 
                           n10538, ZN => n1707);
   U8390 : OAI22_X1 port map( A1 => n11300, A2 => n11538, B1 => n8867, B2 => 
                           n10538, ZN => n1708);
   U8391 : OAI22_X1 port map( A1 => n11300, A2 => n11542, B1 => n8866, B2 => 
                           n11408, ZN => n1709);
   U8392 : OAI22_X1 port map( A1 => n11300, A2 => n11546, B1 => n8865, B2 => 
                           n11408, ZN => n1710);
   U8393 : OAI22_X1 port map( A1 => n11300, A2 => n11550, B1 => n8864, B2 => 
                           n11408, ZN => n1711);
   U8394 : OAI22_X1 port map( A1 => n11300, A2 => n11554, B1 => n8863, B2 => 
                           n11408, ZN => n1712);
   U8395 : OAI22_X1 port map( A1 => n11300, A2 => n11558, B1 => n8862, B2 => 
                           n11408, ZN => n1713);
   U8396 : OAI22_X1 port map( A1 => n11299, A2 => n11562, B1 => n8861, B2 => 
                           n11408, ZN => n1714);
   U8397 : OAI22_X1 port map( A1 => n11299, A2 => n11566, B1 => n8860, B2 => 
                           n11408, ZN => n1715);
   U8398 : OAI22_X1 port map( A1 => n11299, A2 => n11570, B1 => n8859, B2 => 
                           n11408, ZN => n1716);
   U8399 : OAI22_X1 port map( A1 => n11299, A2 => n11574, B1 => n8858, B2 => 
                           n11408, ZN => n1717);
   U8400 : OAI22_X1 port map( A1 => n11299, A2 => n11578, B1 => n8857, B2 => 
                           n10538, ZN => n1718);
   U8401 : OAI22_X1 port map( A1 => n11299, A2 => n11582, B1 => n8856, B2 => 
                           n10538, ZN => n1719);
   U8402 : OAI22_X1 port map( A1 => n11299, A2 => n11586, B1 => n8855, B2 => 
                           n10538, ZN => n1720);
   U8403 : OAI22_X1 port map( A1 => n11299, A2 => n11590, B1 => n8854, B2 => 
                           n10538, ZN => n1721);
   U8404 : OAI22_X1 port map( A1 => n11299, A2 => n11594, B1 => n8853, B2 => 
                           n10538, ZN => n1722);
   U8405 : OAI22_X1 port map( A1 => n11299, A2 => n11598, B1 => n8852, B2 => 
                           n10538, ZN => n1723);
   U8406 : OAI22_X1 port map( A1 => n11299, A2 => n11602, B1 => n8851, B2 => 
                           n10538, ZN => n1724);
   U8407 : OAI22_X1 port map( A1 => n11299, A2 => n11610, B1 => n8850, B2 => 
                           n10538, ZN => n1725);
   U8408 : OAI22_X1 port map( A1 => n11307, A2 => n11482, B1 => n8817, B2 => 
                           n11416, ZN => n1758);
   U8409 : OAI22_X1 port map( A1 => n11307, A2 => n11486, B1 => n8816, B2 => 
                           n11416, ZN => n1759);
   U8410 : OAI22_X1 port map( A1 => n11307, A2 => n11490, B1 => n8815, B2 => 
                           n11416, ZN => n1760);
   U8411 : OAI22_X1 port map( A1 => n11307, A2 => n11494, B1 => n8814, B2 => 
                           n11416, ZN => n1761);
   U8412 : OAI22_X1 port map( A1 => n11307, A2 => n11498, B1 => n8813, B2 => 
                           n11416, ZN => n1762);
   U8413 : OAI22_X1 port map( A1 => n11307, A2 => n11502, B1 => n8812, B2 => 
                           n11416, ZN => n1763);
   U8414 : OAI22_X1 port map( A1 => n11307, A2 => n11506, B1 => n8811, B2 => 
                           n11416, ZN => n1764);
   U8415 : OAI22_X1 port map( A1 => n11307, A2 => n11510, B1 => n8810, B2 => 
                           n11416, ZN => n1765);
   U8416 : OAI22_X1 port map( A1 => n11306, A2 => n11514, B1 => n8809, B2 => 
                           n11416, ZN => n1766);
   U8417 : OAI22_X1 port map( A1 => n11306, A2 => n11518, B1 => n8808, B2 => 
                           n11416, ZN => n1767);
   U8418 : OAI22_X1 port map( A1 => n11306, A2 => n11522, B1 => n8807, B2 => 
                           n11416, ZN => n1768);
   U8419 : OAI22_X1 port map( A1 => n11306, A2 => n11526, B1 => n8806, B2 => 
                           n11416, ZN => n1769);
   U8420 : OAI22_X1 port map( A1 => n11306, A2 => n11530, B1 => n8805, B2 => 
                           n10535, ZN => n1770);
   U8421 : OAI22_X1 port map( A1 => n11306, A2 => n11534, B1 => n8804, B2 => 
                           n10535, ZN => n1771);
   U8422 : OAI22_X1 port map( A1 => n11306, A2 => n11538, B1 => n8803, B2 => 
                           n10535, ZN => n1772);
   U8423 : OAI22_X1 port map( A1 => n11306, A2 => n11542, B1 => n8802, B2 => 
                           n11416, ZN => n1773);
   U8424 : OAI22_X1 port map( A1 => n11306, A2 => n11546, B1 => n8801, B2 => 
                           n11416, ZN => n1774);
   U8425 : OAI22_X1 port map( A1 => n11306, A2 => n11550, B1 => n8800, B2 => 
                           n11416, ZN => n1775);
   U8426 : OAI22_X1 port map( A1 => n11306, A2 => n11554, B1 => n8799, B2 => 
                           n11416, ZN => n1776);
   U8427 : OAI22_X1 port map( A1 => n11306, A2 => n11558, B1 => n8798, B2 => 
                           n11416, ZN => n1777);
   U8428 : OAI22_X1 port map( A1 => n11305, A2 => n11562, B1 => n8797, B2 => 
                           n11416, ZN => n1778);
   U8429 : OAI22_X1 port map( A1 => n11305, A2 => n11566, B1 => n8796, B2 => 
                           n11416, ZN => n1779);
   U8430 : OAI22_X1 port map( A1 => n11305, A2 => n11570, B1 => n8795, B2 => 
                           n11416, ZN => n1780);
   U8431 : OAI22_X1 port map( A1 => n11305, A2 => n11574, B1 => n8794, B2 => 
                           n11416, ZN => n1781);
   U8432 : OAI22_X1 port map( A1 => n11305, A2 => n11578, B1 => n8793, B2 => 
                           n10535, ZN => n1782);
   U8433 : OAI22_X1 port map( A1 => n11305, A2 => n11582, B1 => n8792, B2 => 
                           n10535, ZN => n1783);
   U8434 : OAI22_X1 port map( A1 => n11305, A2 => n11586, B1 => n8791, B2 => 
                           n10535, ZN => n1784);
   U8435 : OAI22_X1 port map( A1 => n11305, A2 => n11590, B1 => n8790, B2 => 
                           n10535, ZN => n1785);
   U8436 : OAI22_X1 port map( A1 => n11305, A2 => n11594, B1 => n8789, B2 => 
                           n10535, ZN => n1786);
   U8437 : OAI22_X1 port map( A1 => n11305, A2 => n11598, B1 => n8788, B2 => 
                           n10535, ZN => n1787);
   U8438 : OAI22_X1 port map( A1 => n11305, A2 => n11602, B1 => n8787, B2 => 
                           n10535, ZN => n1788);
   U8439 : OAI22_X1 port map( A1 => n11305, A2 => n11610, B1 => n8786, B2 => 
                           n10535, ZN => n1789);
   U8440 : OAI22_X1 port map( A1 => n11343, A2 => n11481, B1 => n8433, B2 => 
                           n11464, ZN => n2142);
   U8441 : OAI22_X1 port map( A1 => n11343, A2 => n11485, B1 => n8432, B2 => 
                           n11464, ZN => n2143);
   U8442 : OAI22_X1 port map( A1 => n11343, A2 => n11489, B1 => n8431, B2 => 
                           n11464, ZN => n2144);
   U8443 : OAI22_X1 port map( A1 => n11343, A2 => n11493, B1 => n8430, B2 => 
                           n11464, ZN => n2145);
   U8444 : OAI22_X1 port map( A1 => n11343, A2 => n11497, B1 => n8429, B2 => 
                           n11464, ZN => n2146);
   U8445 : OAI22_X1 port map( A1 => n11343, A2 => n11501, B1 => n8428, B2 => 
                           n11464, ZN => n2147);
   U8446 : OAI22_X1 port map( A1 => n11343, A2 => n11505, B1 => n8427, B2 => 
                           n11464, ZN => n2148);
   U8447 : OAI22_X1 port map( A1 => n11343, A2 => n11509, B1 => n8426, B2 => 
                           n11464, ZN => n2149);
   U8448 : OAI22_X1 port map( A1 => n11342, A2 => n11513, B1 => n8425, B2 => 
                           n11464, ZN => n2150);
   U8449 : OAI22_X1 port map( A1 => n11342, A2 => n11517, B1 => n8424, B2 => 
                           n11464, ZN => n2151);
   U8450 : OAI22_X1 port map( A1 => n11342, A2 => n11521, B1 => n8423, B2 => 
                           n11464, ZN => n2152);
   U8451 : OAI22_X1 port map( A1 => n11342, A2 => n11525, B1 => n8422, B2 => 
                           n11464, ZN => n2153);
   U8452 : OAI22_X1 port map( A1 => n11342, A2 => n11529, B1 => n8421, B2 => 
                           n10520, ZN => n2154);
   U8453 : OAI22_X1 port map( A1 => n11342, A2 => n11533, B1 => n8420, B2 => 
                           n10520, ZN => n2155);
   U8454 : OAI22_X1 port map( A1 => n11342, A2 => n11537, B1 => n8419, B2 => 
                           n10520, ZN => n2156);
   U8455 : OAI22_X1 port map( A1 => n11342, A2 => n11541, B1 => n8418, B2 => 
                           n11464, ZN => n2157);
   U8456 : OAI22_X1 port map( A1 => n11342, A2 => n11545, B1 => n8417, B2 => 
                           n11464, ZN => n2158);
   U8457 : OAI22_X1 port map( A1 => n11342, A2 => n11549, B1 => n8416, B2 => 
                           n11464, ZN => n2159);
   U8458 : OAI22_X1 port map( A1 => n11342, A2 => n11553, B1 => n8415, B2 => 
                           n11464, ZN => n2160);
   U8459 : OAI22_X1 port map( A1 => n11342, A2 => n11557, B1 => n8414, B2 => 
                           n11464, ZN => n2161);
   U8460 : OAI22_X1 port map( A1 => n11341, A2 => n11561, B1 => n8413, B2 => 
                           n11464, ZN => n2162);
   U8461 : OAI22_X1 port map( A1 => n11341, A2 => n11565, B1 => n8412, B2 => 
                           n11464, ZN => n2163);
   U8462 : OAI22_X1 port map( A1 => n11341, A2 => n11569, B1 => n8411, B2 => 
                           n11464, ZN => n2164);
   U8463 : OAI22_X1 port map( A1 => n11341, A2 => n11573, B1 => n8410, B2 => 
                           n11464, ZN => n2165);
   U8464 : OAI22_X1 port map( A1 => n11341, A2 => n11577, B1 => n8409, B2 => 
                           n10520, ZN => n2166);
   U8465 : OAI22_X1 port map( A1 => n11341, A2 => n11581, B1 => n8408, B2 => 
                           n10520, ZN => n2167);
   U8466 : OAI22_X1 port map( A1 => n11341, A2 => n11585, B1 => n8407, B2 => 
                           n10520, ZN => n2168);
   U8467 : OAI22_X1 port map( A1 => n11341, A2 => n11589, B1 => n8406, B2 => 
                           n10520, ZN => n2169);
   U8468 : OAI22_X1 port map( A1 => n11341, A2 => n11593, B1 => n8405, B2 => 
                           n10520, ZN => n2170);
   U8469 : OAI22_X1 port map( A1 => n11341, A2 => n11597, B1 => n8404, B2 => 
                           n10520, ZN => n2171);
   U8470 : OAI22_X1 port map( A1 => n11341, A2 => n11601, B1 => n8403, B2 => 
                           n10520, ZN => n2172);
   U8471 : OAI22_X1 port map( A1 => n11341, A2 => n11609, B1 => n8402, B2 => 
                           n10520, ZN => n2173);
   U8472 : OAI22_X1 port map( A1 => n11316, A2 => n11482, B1 => n8721, B2 => 
                           n11428, ZN => n1854);
   U8473 : OAI22_X1 port map( A1 => n11316, A2 => n11486, B1 => n8720, B2 => 
                           n11428, ZN => n1855);
   U8474 : OAI22_X1 port map( A1 => n11316, A2 => n11490, B1 => n8719, B2 => 
                           n11428, ZN => n1856);
   U8475 : OAI22_X1 port map( A1 => n11316, A2 => n11494, B1 => n8718, B2 => 
                           n11428, ZN => n1857);
   U8476 : OAI22_X1 port map( A1 => n11316, A2 => n11498, B1 => n8717, B2 => 
                           n11428, ZN => n1858);
   U8477 : OAI22_X1 port map( A1 => n11316, A2 => n11502, B1 => n8716, B2 => 
                           n11428, ZN => n1859);
   U8478 : OAI22_X1 port map( A1 => n11316, A2 => n11506, B1 => n8715, B2 => 
                           n11428, ZN => n1860);
   U8479 : OAI22_X1 port map( A1 => n11316, A2 => n11510, B1 => n8714, B2 => 
                           n11428, ZN => n1861);
   U8480 : OAI22_X1 port map( A1 => n11315, A2 => n11514, B1 => n8713, B2 => 
                           n11428, ZN => n1862);
   U8481 : OAI22_X1 port map( A1 => n11315, A2 => n11518, B1 => n8712, B2 => 
                           n11428, ZN => n1863);
   U8482 : OAI22_X1 port map( A1 => n11315, A2 => n11522, B1 => n8711, B2 => 
                           n11428, ZN => n1864);
   U8483 : OAI22_X1 port map( A1 => n11315, A2 => n11526, B1 => n8710, B2 => 
                           n11428, ZN => n1865);
   U8484 : OAI22_X1 port map( A1 => n11315, A2 => n11530, B1 => n8709, B2 => 
                           n10532, ZN => n1866);
   U8485 : OAI22_X1 port map( A1 => n11315, A2 => n11534, B1 => n8708, B2 => 
                           n10532, ZN => n1867);
   U8486 : OAI22_X1 port map( A1 => n11315, A2 => n11538, B1 => n8707, B2 => 
                           n10532, ZN => n1868);
   U8487 : OAI22_X1 port map( A1 => n11315, A2 => n11542, B1 => n8706, B2 => 
                           n11428, ZN => n1869);
   U8488 : OAI22_X1 port map( A1 => n11315, A2 => n11546, B1 => n8705, B2 => 
                           n11428, ZN => n1870);
   U8489 : OAI22_X1 port map( A1 => n11315, A2 => n11550, B1 => n8704, B2 => 
                           n11428, ZN => n1871);
   U8490 : OAI22_X1 port map( A1 => n11315, A2 => n11554, B1 => n8703, B2 => 
                           n11428, ZN => n1872);
   U8491 : OAI22_X1 port map( A1 => n11315, A2 => n11558, B1 => n8702, B2 => 
                           n11428, ZN => n1873);
   U8492 : OAI22_X1 port map( A1 => n11314, A2 => n11562, B1 => n8701, B2 => 
                           n11428, ZN => n1874);
   U8493 : OAI22_X1 port map( A1 => n11314, A2 => n11566, B1 => n8700, B2 => 
                           n11428, ZN => n1875);
   U8494 : OAI22_X1 port map( A1 => n11314, A2 => n11570, B1 => n8699, B2 => 
                           n11428, ZN => n1876);
   U8495 : OAI22_X1 port map( A1 => n11314, A2 => n11574, B1 => n8698, B2 => 
                           n11428, ZN => n1877);
   U8496 : OAI22_X1 port map( A1 => n11314, A2 => n11578, B1 => n8697, B2 => 
                           n10532, ZN => n1878);
   U8497 : OAI22_X1 port map( A1 => n11314, A2 => n11582, B1 => n8696, B2 => 
                           n10532, ZN => n1879);
   U8498 : OAI22_X1 port map( A1 => n11314, A2 => n11586, B1 => n8695, B2 => 
                           n10532, ZN => n1880);
   U8499 : OAI22_X1 port map( A1 => n11314, A2 => n11590, B1 => n8694, B2 => 
                           n10532, ZN => n1881);
   U8500 : OAI22_X1 port map( A1 => n11314, A2 => n11594, B1 => n8693, B2 => 
                           n10532, ZN => n1882);
   U8501 : OAI22_X1 port map( A1 => n11314, A2 => n11598, B1 => n8692, B2 => 
                           n10532, ZN => n1883);
   U8502 : OAI22_X1 port map( A1 => n11314, A2 => n11602, B1 => n8691, B2 => 
                           n10532, ZN => n1884);
   U8503 : OAI22_X1 port map( A1 => n11314, A2 => n11610, B1 => n8690, B2 => 
                           n10532, ZN => n1885);
   U8504 : OAI22_X1 port map( A1 => n11349, A2 => n11501, B1 => n8364, B2 => 
                           n11472, ZN => n2211);
   U8505 : OAI22_X1 port map( A1 => n11349, A2 => n11505, B1 => n8363, B2 => 
                           n11472, ZN => n2212);
   U8506 : OAI22_X1 port map( A1 => n11349, A2 => n11509, B1 => n8362, B2 => 
                           n11472, ZN => n2213);
   U8507 : OAI22_X1 port map( A1 => n11348, A2 => n11517, B1 => n8360, B2 => 
                           n11472, ZN => n2215);
   U8508 : OAI22_X1 port map( A1 => n11348, A2 => n11521, B1 => n8359, B2 => 
                           n11472, ZN => n2216);
   U8509 : OAI22_X1 port map( A1 => n11348, A2 => n11525, B1 => n8358, B2 => 
                           n11472, ZN => n2217);
   U8510 : OAI22_X1 port map( A1 => n11348, A2 => n11529, B1 => n8357, B2 => 
                           n10515, ZN => n2218);
   U8511 : OAI22_X1 port map( A1 => n11348, A2 => n11533, B1 => n8356, B2 => 
                           n10515, ZN => n2219);
   U8512 : OAI22_X1 port map( A1 => n11348, A2 => n11541, B1 => n8354, B2 => 
                           n10515, ZN => n2221);
   U8513 : OAI22_X1 port map( A1 => n11348, A2 => n11549, B1 => n8352, B2 => 
                           n11472, ZN => n2223);
   U8514 : OAI22_X1 port map( A1 => n11348, A2 => n11553, B1 => n8351, B2 => 
                           n11472, ZN => n2224);
   U8515 : OAI22_X1 port map( A1 => n11347, A2 => n11561, B1 => n8349, B2 => 
                           n11472, ZN => n2226);
   U8516 : OAI22_X1 port map( A1 => n11347, A2 => n11573, B1 => n8346, B2 => 
                           n11472, ZN => n2229);
   U8517 : OAI22_X1 port map( A1 => n11347, A2 => n11589, B1 => n8342, B2 => 
                           n10515, ZN => n2233);
   U8518 : OAI22_X1 port map( A1 => n11347, A2 => n11593, B1 => n8341, B2 => 
                           n10515, ZN => n2234);
   U8519 : OAI22_X1 port map( A1 => n11347, A2 => n11609, B1 => n8338, B2 => 
                           n10515, ZN => n2237);
   U8520 : OAI22_X1 port map( A1 => n11264, A2 => n11515, B1 => n9257, B2 => 
                           n11360, ZN => n1318);
   U8521 : OAI22_X1 port map( A1 => n11264, A2 => n11519, B1 => n9256, B2 => 
                           n11360, ZN => n1319);
   U8522 : OAI22_X1 port map( A1 => n11264, A2 => n11523, B1 => n9255, B2 => 
                           n11360, ZN => n1320);
   U8523 : OAI22_X1 port map( A1 => n11264, A2 => n11527, B1 => n9254, B2 => 
                           n11360, ZN => n1321);
   U8524 : OAI22_X1 port map( A1 => n11264, A2 => n11531, B1 => n9253, B2 => 
                           n10554, ZN => n1322);
   U8525 : OAI22_X1 port map( A1 => n11264, A2 => n11535, B1 => n9252, B2 => 
                           n10554, ZN => n1323);
   U8526 : OAI22_X1 port map( A1 => n11264, A2 => n11539, B1 => n9251, B2 => 
                           n10554, ZN => n1324);
   U8527 : OAI22_X1 port map( A1 => n11264, A2 => n11543, B1 => n9250, B2 => 
                           n11360, ZN => n1325);
   U8528 : OAI22_X1 port map( A1 => n11264, A2 => n11547, B1 => n9249, B2 => 
                           n11360, ZN => n1326);
   U8529 : OAI22_X1 port map( A1 => n11264, A2 => n11551, B1 => n9248, B2 => 
                           n11360, ZN => n1327);
   U8530 : OAI22_X1 port map( A1 => n11264, A2 => n11555, B1 => n9247, B2 => 
                           n11360, ZN => n1328);
   U8531 : OAI22_X1 port map( A1 => n11264, A2 => n11559, B1 => n9246, B2 => 
                           n11360, ZN => n1329);
   U8532 : OAI22_X1 port map( A1 => n11263, A2 => n11567, B1 => n9244, B2 => 
                           n11360, ZN => n1331);
   U8533 : OAI22_X1 port map( A1 => n11263, A2 => n11571, B1 => n9243, B2 => 
                           n11360, ZN => n1332);
   U8534 : OAI22_X1 port map( A1 => n11263, A2 => n11575, B1 => n9242, B2 => 
                           n11360, ZN => n1333);
   U8535 : OAI22_X1 port map( A1 => n11263, A2 => n11579, B1 => n9241, B2 => 
                           n10554, ZN => n1334);
   U8536 : OAI22_X1 port map( A1 => n11263, A2 => n11583, B1 => n9240, B2 => 
                           n10554, ZN => n1335);
   U8537 : OAI22_X1 port map( A1 => n11263, A2 => n11591, B1 => n9238, B2 => 
                           n10554, ZN => n1337);
   U8538 : OAI22_X1 port map( A1 => n11263, A2 => n11599, B1 => n9236, B2 => 
                           n10554, ZN => n1339);
   U8539 : OAI22_X1 port map( A1 => n11263, A2 => n11603, B1 => n9235, B2 => 
                           n10554, ZN => n1340);
   U8540 : OAI22_X1 port map( A1 => n11263, A2 => n11611, B1 => n9234, B2 => 
                           n10554, ZN => n1341);
   U8541 : OAI22_X1 port map( A1 => n11280, A2 => n11483, B1 => n9105, B2 => 
                           n11380, ZN => n1470);
   U8542 : OAI22_X1 port map( A1 => n11280, A2 => n11491, B1 => n9103, B2 => 
                           n11380, ZN => n1472);
   U8543 : OAI22_X1 port map( A1 => n11280, A2 => n11503, B1 => n9100, B2 => 
                           n11380, ZN => n1475);
   U8544 : OAI22_X1 port map( A1 => n11280, A2 => n11507, B1 => n9099, B2 => 
                           n11380, ZN => n1476);
   U8545 : OAI22_X1 port map( A1 => n11280, A2 => n11511, B1 => n9098, B2 => 
                           n11380, ZN => n1477);
   U8546 : OAI22_X1 port map( A1 => n11279, A2 => n11515, B1 => n9097, B2 => 
                           n11380, ZN => n1478);
   U8547 : OAI22_X1 port map( A1 => n11279, A2 => n11519, B1 => n9096, B2 => 
                           n11380, ZN => n1479);
   U8548 : OAI22_X1 port map( A1 => n11279, A2 => n11523, B1 => n9095, B2 => 
                           n11380, ZN => n1480);
   U8549 : OAI22_X1 port map( A1 => n11279, A2 => n11527, B1 => n9094, B2 => 
                           n11380, ZN => n1481);
   U8550 : OAI22_X1 port map( A1 => n11279, A2 => n11543, B1 => n9090, B2 => 
                           n10548, ZN => n1485);
   U8551 : OAI22_X1 port map( A1 => n11279, A2 => n11547, B1 => n9089, B2 => 
                           n10548, ZN => n1486);
   U8552 : OAI22_X1 port map( A1 => n11279, A2 => n11551, B1 => n9088, B2 => 
                           n10548, ZN => n1487);
   U8553 : OAI22_X1 port map( A1 => n11279, A2 => n11559, B1 => n9086, B2 => 
                           n11380, ZN => n1489);
   U8554 : OAI22_X1 port map( A1 => n11278, A2 => n11563, B1 => n9085, B2 => 
                           n11380, ZN => n1490);
   U8555 : OAI22_X1 port map( A1 => n11278, A2 => n11567, B1 => n9084, B2 => 
                           n11380, ZN => n1491);
   U8556 : OAI22_X1 port map( A1 => n11278, A2 => n11571, B1 => n9083, B2 => 
                           n11380, ZN => n1492);
   U8557 : OAI22_X1 port map( A1 => n11278, A2 => n11575, B1 => n9082, B2 => 
                           n11380, ZN => n1493);
   U8558 : OAI22_X1 port map( A1 => n11278, A2 => n11579, B1 => n9081, B2 => 
                           n10548, ZN => n1494);
   U8559 : OAI22_X1 port map( A1 => n11278, A2 => n11587, B1 => n9079, B2 => 
                           n10548, ZN => n1496);
   U8560 : OAI22_X1 port map( A1 => n11278, A2 => n11591, B1 => n9078, B2 => 
                           n10548, ZN => n1497);
   U8561 : OAI22_X1 port map( A1 => n11278, A2 => n11595, B1 => n9077, B2 => 
                           n10548, ZN => n1498);
   U8562 : OAI22_X1 port map( A1 => n11278, A2 => n11599, B1 => n9076, B2 => 
                           n10548, ZN => n1499);
   U8563 : OAI22_X1 port map( A1 => n11278, A2 => n11611, B1 => n9074, B2 => 
                           n10548, ZN => n1501);
   U8564 : OAI22_X1 port map( A1 => n11292, A2 => n11482, B1 => n8977, B2 => 
                           n11396, ZN => n1598);
   U8565 : OAI22_X1 port map( A1 => n11292, A2 => n11486, B1 => n8976, B2 => 
                           n11396, ZN => n1599);
   U8566 : OAI22_X1 port map( A1 => n11292, A2 => n11490, B1 => n8975, B2 => 
                           n11396, ZN => n1600);
   U8567 : OAI22_X1 port map( A1 => n11292, A2 => n11494, B1 => n8974, B2 => 
                           n11396, ZN => n1601);
   U8568 : OAI22_X1 port map( A1 => n11292, A2 => n11502, B1 => n8972, B2 => 
                           n11396, ZN => n1603);
   U8569 : OAI22_X1 port map( A1 => n11292, A2 => n11506, B1 => n8971, B2 => 
                           n11396, ZN => n1604);
   U8570 : OAI22_X1 port map( A1 => n11292, A2 => n11510, B1 => n8970, B2 => 
                           n11396, ZN => n1605);
   U8571 : OAI22_X1 port map( A1 => n11291, A2 => n11514, B1 => n8969, B2 => 
                           n11396, ZN => n1606);
   U8572 : OAI22_X1 port map( A1 => n11291, A2 => n11522, B1 => n8967, B2 => 
                           n11396, ZN => n1608);
   U8573 : OAI22_X1 port map( A1 => n11291, A2 => n11526, B1 => n8966, B2 => 
                           n11396, ZN => n1609);
   U8574 : OAI22_X1 port map( A1 => n11291, A2 => n11530, B1 => n8965, B2 => 
                           n10543, ZN => n1610);
   U8575 : OAI22_X1 port map( A1 => n11291, A2 => n11534, B1 => n8964, B2 => 
                           n10543, ZN => n1611);
   U8576 : OAI22_X1 port map( A1 => n11291, A2 => n11538, B1 => n8963, B2 => 
                           n10543, ZN => n1612);
   U8577 : OAI22_X1 port map( A1 => n11291, A2 => n11542, B1 => n8962, B2 => 
                           n11396, ZN => n1613);
   U8578 : OAI22_X1 port map( A1 => n11291, A2 => n11546, B1 => n8961, B2 => 
                           n11396, ZN => n1614);
   U8579 : OAI22_X1 port map( A1 => n11291, A2 => n11550, B1 => n8960, B2 => 
                           n11396, ZN => n1615);
   U8580 : OAI22_X1 port map( A1 => n11291, A2 => n11554, B1 => n8959, B2 => 
                           n11396, ZN => n1616);
   U8581 : OAI22_X1 port map( A1 => n11291, A2 => n11558, B1 => n8958, B2 => 
                           n11396, ZN => n1617);
   U8582 : OAI22_X1 port map( A1 => n11290, A2 => n11562, B1 => n8957, B2 => 
                           n11396, ZN => n1618);
   U8583 : OAI22_X1 port map( A1 => n11290, A2 => n11570, B1 => n8955, B2 => 
                           n11396, ZN => n1620);
   U8584 : OAI22_X1 port map( A1 => n11290, A2 => n11574, B1 => n8954, B2 => 
                           n11396, ZN => n1621);
   U8585 : OAI22_X1 port map( A1 => n11290, A2 => n11578, B1 => n8953, B2 => 
                           n10543, ZN => n1622);
   U8586 : OAI22_X1 port map( A1 => n11290, A2 => n11582, B1 => n8952, B2 => 
                           n10543, ZN => n1623);
   U8587 : OAI22_X1 port map( A1 => n11290, A2 => n11586, B1 => n8951, B2 => 
                           n10543, ZN => n1624);
   U8588 : OAI22_X1 port map( A1 => n11290, A2 => n11590, B1 => n8950, B2 => 
                           n10543, ZN => n1625);
   U8589 : OAI22_X1 port map( A1 => n11290, A2 => n11594, B1 => n8949, B2 => 
                           n10543, ZN => n1626);
   U8590 : OAI22_X1 port map( A1 => n11290, A2 => n11598, B1 => n8948, B2 => 
                           n10543, ZN => n1627);
   U8591 : OAI22_X1 port map( A1 => n11290, A2 => n11602, B1 => n8947, B2 => 
                           n10543, ZN => n1628);
   U8592 : OAI22_X1 port map( A1 => n11295, A2 => n11482, B1 => n8945, B2 => 
                           n11400, ZN => n1630);
   U8593 : OAI22_X1 port map( A1 => n11295, A2 => n11486, B1 => n8944, B2 => 
                           n11400, ZN => n1631);
   U8594 : OAI22_X1 port map( A1 => n11295, A2 => n11490, B1 => n8943, B2 => 
                           n11400, ZN => n1632);
   U8595 : OAI22_X1 port map( A1 => n11295, A2 => n11494, B1 => n8942, B2 => 
                           n11400, ZN => n1633);
   U8596 : OAI22_X1 port map( A1 => n11295, A2 => n11498, B1 => n8941, B2 => 
                           n11400, ZN => n1634);
   U8597 : OAI22_X1 port map( A1 => n11295, A2 => n11506, B1 => n8939, B2 => 
                           n11400, ZN => n1636);
   U8598 : OAI22_X1 port map( A1 => n11295, A2 => n11510, B1 => n8938, B2 => 
                           n11400, ZN => n1637);
   U8599 : OAI22_X1 port map( A1 => n11294, A2 => n11514, B1 => n8937, B2 => 
                           n11400, ZN => n1638);
   U8600 : OAI22_X1 port map( A1 => n11294, A2 => n11518, B1 => n8936, B2 => 
                           n11400, ZN => n1639);
   U8601 : OAI22_X1 port map( A1 => n11294, A2 => n11522, B1 => n8935, B2 => 
                           n11400, ZN => n1640);
   U8602 : OAI22_X1 port map( A1 => n11294, A2 => n11526, B1 => n8934, B2 => 
                           n11400, ZN => n1641);
   U8603 : OAI22_X1 port map( A1 => n11294, A2 => n11530, B1 => n8933, B2 => 
                           n10541, ZN => n1642);
   U8604 : OAI22_X1 port map( A1 => n11294, A2 => n11534, B1 => n8932, B2 => 
                           n10541, ZN => n1643);
   U8605 : OAI22_X1 port map( A1 => n11294, A2 => n11538, B1 => n8931, B2 => 
                           n10541, ZN => n1644);
   U8606 : OAI22_X1 port map( A1 => n11294, A2 => n11542, B1 => n8930, B2 => 
                           n11400, ZN => n1645);
   U8607 : OAI22_X1 port map( A1 => n11294, A2 => n11546, B1 => n8929, B2 => 
                           n11400, ZN => n1646);
   U8608 : OAI22_X1 port map( A1 => n11294, A2 => n11554, B1 => n8927, B2 => 
                           n11400, ZN => n1648);
   U8609 : OAI22_X1 port map( A1 => n11294, A2 => n11558, B1 => n8926, B2 => 
                           n11400, ZN => n1649);
   U8610 : OAI22_X1 port map( A1 => n11293, A2 => n11562, B1 => n8925, B2 => 
                           n11400, ZN => n1650);
   U8611 : OAI22_X1 port map( A1 => n11293, A2 => n11570, B1 => n8923, B2 => 
                           n11400, ZN => n1652);
   U8612 : OAI22_X1 port map( A1 => n11293, A2 => n11574, B1 => n8922, B2 => 
                           n11400, ZN => n1653);
   U8613 : OAI22_X1 port map( A1 => n11293, A2 => n11578, B1 => n8921, B2 => 
                           n10541, ZN => n1654);
   U8614 : OAI22_X1 port map( A1 => n11293, A2 => n11582, B1 => n8920, B2 => 
                           n10541, ZN => n1655);
   U8615 : OAI22_X1 port map( A1 => n11293, A2 => n11586, B1 => n8919, B2 => 
                           n10541, ZN => n1656);
   U8616 : OAI22_X1 port map( A1 => n11293, A2 => n11590, B1 => n8918, B2 => 
                           n10541, ZN => n1657);
   U8617 : OAI22_X1 port map( A1 => n11293, A2 => n11594, B1 => n8917, B2 => 
                           n10541, ZN => n1658);
   U8618 : OAI22_X1 port map( A1 => n11293, A2 => n11598, B1 => n8916, B2 => 
                           n10541, ZN => n1659);
   U8619 : OAI22_X1 port map( A1 => n11293, A2 => n11610, B1 => n8914, B2 => 
                           n10541, ZN => n1661);
   U8620 : OAI22_X1 port map( A1 => n11319, A2 => n11490, B1 => n8687, B2 => 
                           n11432, ZN => n1888);
   U8621 : OAI22_X1 port map( A1 => n11319, A2 => n11494, B1 => n8686, B2 => 
                           n11432, ZN => n1889);
   U8622 : OAI22_X1 port map( A1 => n11319, A2 => n11498, B1 => n8685, B2 => 
                           n11432, ZN => n1890);
   U8623 : OAI22_X1 port map( A1 => n11319, A2 => n11502, B1 => n8684, B2 => 
                           n11432, ZN => n1891);
   U8624 : OAI22_X1 port map( A1 => n11319, A2 => n11506, B1 => n8683, B2 => 
                           n11432, ZN => n1892);
   U8625 : OAI22_X1 port map( A1 => n11319, A2 => n11510, B1 => n8682, B2 => 
                           n11432, ZN => n1893);
   U8626 : OAI22_X1 port map( A1 => n11318, A2 => n11514, B1 => n8681, B2 => 
                           n11432, ZN => n1894);
   U8627 : OAI22_X1 port map( A1 => n11318, A2 => n11518, B1 => n8680, B2 => 
                           n11432, ZN => n1895);
   U8628 : OAI22_X1 port map( A1 => n11318, A2 => n11522, B1 => n8679, B2 => 
                           n11432, ZN => n1896);
   U8629 : OAI22_X1 port map( A1 => n11318, A2 => n11526, B1 => n8678, B2 => 
                           n11432, ZN => n1897);
   U8630 : OAI22_X1 port map( A1 => n11318, A2 => n11530, B1 => n8677, B2 => 
                           n10530, ZN => n1898);
   U8631 : OAI22_X1 port map( A1 => n11318, A2 => n11534, B1 => n8676, B2 => 
                           n10530, ZN => n1899);
   U8632 : OAI22_X1 port map( A1 => n11318, A2 => n11542, B1 => n8674, B2 => 
                           n10530, ZN => n1901);
   U8633 : OAI22_X1 port map( A1 => n11318, A2 => n11546, B1 => n8673, B2 => 
                           n11432, ZN => n1902);
   U8634 : OAI22_X1 port map( A1 => n11318, A2 => n11550, B1 => n8672, B2 => 
                           n11432, ZN => n1903);
   U8635 : OAI22_X1 port map( A1 => n11318, A2 => n11554, B1 => n8671, B2 => 
                           n11432, ZN => n1904);
   U8636 : OAI22_X1 port map( A1 => n11317, A2 => n11566, B1 => n8668, B2 => 
                           n11432, ZN => n1907);
   U8637 : OAI22_X1 port map( A1 => n11317, A2 => n11574, B1 => n8666, B2 => 
                           n11432, ZN => n1909);
   U8638 : OAI22_X1 port map( A1 => n11317, A2 => n11578, B1 => n8665, B2 => 
                           n10530, ZN => n1910);
   U8639 : OAI22_X1 port map( A1 => n11317, A2 => n11582, B1 => n8664, B2 => 
                           n10530, ZN => n1911);
   U8640 : OAI22_X1 port map( A1 => n11317, A2 => n11586, B1 => n8663, B2 => 
                           n10530, ZN => n1912);
   U8641 : OAI22_X1 port map( A1 => n11317, A2 => n11590, B1 => n8662, B2 => 
                           n10530, ZN => n1913);
   U8642 : OAI22_X1 port map( A1 => n11317, A2 => n11594, B1 => n8661, B2 => 
                           n10530, ZN => n1914);
   U8643 : OAI22_X1 port map( A1 => n11317, A2 => n11598, B1 => n8660, B2 => 
                           n10530, ZN => n1915);
   U8644 : OAI22_X1 port map( A1 => n11317, A2 => n11602, B1 => n8659, B2 => 
                           n10530, ZN => n1916);
   U8645 : OAI22_X1 port map( A1 => n11317, A2 => n11610, B1 => n8658, B2 => 
                           n10530, ZN => n1917);
   U8646 : OAI22_X1 port map( A1 => n11349, A2 => n11481, B1 => n8369, B2 => 
                           n11472, ZN => n2206);
   U8647 : OAI22_X1 port map( A1 => n11349, A2 => n11485, B1 => n8368, B2 => 
                           n11472, ZN => n2207);
   U8648 : OAI22_X1 port map( A1 => n11349, A2 => n11489, B1 => n8367, B2 => 
                           n11472, ZN => n2208);
   U8649 : OAI22_X1 port map( A1 => n11349, A2 => n11493, B1 => n8366, B2 => 
                           n11472, ZN => n2209);
   U8650 : OAI22_X1 port map( A1 => n11349, A2 => n11497, B1 => n8365, B2 => 
                           n11472, ZN => n2210);
   U8651 : OAI22_X1 port map( A1 => n11348, A2 => n11537, B1 => n8355, B2 => 
                           n11472, ZN => n2220);
   U8652 : OAI22_X1 port map( A1 => n11348, A2 => n11545, B1 => n8353, B2 => 
                           n11472, ZN => n2222);
   U8653 : OAI22_X1 port map( A1 => n11347, A2 => n11581, B1 => n8344, B2 => 
                           n10515, ZN => n2231);
   U8654 : OAI22_X1 port map( A1 => n11347, A2 => n11597, B1 => n8340, B2 => 
                           n10515, ZN => n2235);
   U8655 : OAI22_X1 port map( A1 => n11347, A2 => n11601, B1 => n8339, B2 => 
                           n10515, ZN => n2236);
   U8656 : OAI22_X1 port map( A1 => n11265, A2 => n11483, B1 => n9265, B2 => 
                           n11360, ZN => n1310);
   U8657 : OAI22_X1 port map( A1 => n11265, A2 => n11487, B1 => n9264, B2 => 
                           n11360, ZN => n1311);
   U8658 : OAI22_X1 port map( A1 => n11265, A2 => n11491, B1 => n9263, B2 => 
                           n11360, ZN => n1312);
   U8659 : OAI22_X1 port map( A1 => n11265, A2 => n11495, B1 => n9262, B2 => 
                           n11360, ZN => n1313);
   U8660 : OAI22_X1 port map( A1 => n11265, A2 => n11499, B1 => n9261, B2 => 
                           n11360, ZN => n1314);
   U8661 : OAI22_X1 port map( A1 => n11265, A2 => n11503, B1 => n9260, B2 => 
                           n11360, ZN => n1315);
   U8662 : OAI22_X1 port map( A1 => n11265, A2 => n11507, B1 => n9259, B2 => 
                           n11360, ZN => n1316);
   U8663 : OAI22_X1 port map( A1 => n11265, A2 => n11511, B1 => n9258, B2 => 
                           n11360, ZN => n1317);
   U8664 : OAI22_X1 port map( A1 => n11263, A2 => n11563, B1 => n9245, B2 => 
                           n11360, ZN => n1330);
   U8665 : OAI22_X1 port map( A1 => n11263, A2 => n11587, B1 => n9239, B2 => 
                           n10554, ZN => n1336);
   U8666 : OAI22_X1 port map( A1 => n11263, A2 => n11595, B1 => n9237, B2 => 
                           n10554, ZN => n1338);
   U8667 : OAI22_X1 port map( A1 => n11280, A2 => n11487, B1 => n9104, B2 => 
                           n11380, ZN => n1471);
   U8668 : OAI22_X1 port map( A1 => n11280, A2 => n11495, B1 => n9102, B2 => 
                           n11380, ZN => n1473);
   U8669 : OAI22_X1 port map( A1 => n11280, A2 => n11499, B1 => n9101, B2 => 
                           n11380, ZN => n1474);
   U8670 : OAI22_X1 port map( A1 => n11279, A2 => n11531, B1 => n9093, B2 => 
                           n11380, ZN => n1482);
   U8671 : OAI22_X1 port map( A1 => n11279, A2 => n11535, B1 => n9092, B2 => 
                           n11380, ZN => n1483);
   U8672 : OAI22_X1 port map( A1 => n11279, A2 => n11539, B1 => n9091, B2 => 
                           n11380, ZN => n1484);
   U8673 : OAI22_X1 port map( A1 => n11279, A2 => n11555, B1 => n9087, B2 => 
                           n11380, ZN => n1488);
   U8674 : OAI22_X1 port map( A1 => n11278, A2 => n11583, B1 => n9080, B2 => 
                           n10548, ZN => n1495);
   U8675 : OAI22_X1 port map( A1 => n11278, A2 => n11603, B1 => n9075, B2 => 
                           n10548, ZN => n1500);
   U8676 : OAI22_X1 port map( A1 => n11292, A2 => n11498, B1 => n8973, B2 => 
                           n11396, ZN => n1602);
   U8677 : OAI22_X1 port map( A1 => n11291, A2 => n11518, B1 => n8968, B2 => 
                           n11396, ZN => n1607);
   U8678 : OAI22_X1 port map( A1 => n11290, A2 => n11566, B1 => n8956, B2 => 
                           n11396, ZN => n1619);
   U8679 : OAI22_X1 port map( A1 => n11290, A2 => n11610, B1 => n8946, B2 => 
                           n10543, ZN => n1629);
   U8680 : OAI22_X1 port map( A1 => n11295, A2 => n11502, B1 => n8940, B2 => 
                           n11400, ZN => n1635);
   U8681 : OAI22_X1 port map( A1 => n11294, A2 => n11550, B1 => n8928, B2 => 
                           n11400, ZN => n1647);
   U8682 : OAI22_X1 port map( A1 => n11293, A2 => n11566, B1 => n8924, B2 => 
                           n11400, ZN => n1651);
   U8683 : OAI22_X1 port map( A1 => n11293, A2 => n11602, B1 => n8915, B2 => 
                           n10541, ZN => n1660);
   U8684 : OAI22_X1 port map( A1 => n11319, A2 => n11482, B1 => n8689, B2 => 
                           n11432, ZN => n1886);
   U8685 : OAI22_X1 port map( A1 => n11319, A2 => n11486, B1 => n8688, B2 => 
                           n11432, ZN => n1887);
   U8686 : OAI22_X1 port map( A1 => n11318, A2 => n11538, B1 => n8675, B2 => 
                           n11432, ZN => n1900);
   U8687 : OAI22_X1 port map( A1 => n11318, A2 => n11558, B1 => n8670, B2 => 
                           n11432, ZN => n1905);
   U8688 : OAI22_X1 port map( A1 => n11317, A2 => n11562, B1 => n8669, B2 => 
                           n11432, ZN => n1906);
   U8689 : OAI22_X1 port map( A1 => n11317, A2 => n11570, B1 => n8667, B2 => 
                           n11432, ZN => n1908);
   U8690 : OAI22_X1 port map( A1 => n11322, A2 => n11481, B1 => n8657, B2 => 
                           n11436, ZN => n1918);
   U8691 : OAI22_X1 port map( A1 => n11322, A2 => n11485, B1 => n8656, B2 => 
                           n11436, ZN => n1919);
   U8692 : OAI22_X1 port map( A1 => n11322, A2 => n11493, B1 => n8654, B2 => 
                           n11436, ZN => n1921);
   U8693 : OAI22_X1 port map( A1 => n11322, A2 => n11497, B1 => n8653, B2 => 
                           n11436, ZN => n1922);
   U8694 : OAI22_X1 port map( A1 => n11322, A2 => n11501, B1 => n8652, B2 => 
                           n11436, ZN => n1923);
   U8695 : OAI22_X1 port map( A1 => n11322, A2 => n11505, B1 => n8651, B2 => 
                           n11436, ZN => n1924);
   U8696 : OAI22_X1 port map( A1 => n11322, A2 => n11509, B1 => n8650, B2 => 
                           n11436, ZN => n1925);
   U8697 : OAI22_X1 port map( A1 => n11321, A2 => n11513, B1 => n8649, B2 => 
                           n11436, ZN => n1926);
   U8698 : OAI22_X1 port map( A1 => n11321, A2 => n11517, B1 => n8648, B2 => 
                           n11436, ZN => n1927);
   U8699 : OAI22_X1 port map( A1 => n11321, A2 => n11521, B1 => n8647, B2 => 
                           n11436, ZN => n1928);
   U8700 : OAI22_X1 port map( A1 => n11321, A2 => n11525, B1 => n8646, B2 => 
                           n11436, ZN => n1929);
   U8701 : OAI22_X1 port map( A1 => n11321, A2 => n11529, B1 => n8645, B2 => 
                           n10529, ZN => n1930);
   U8702 : OAI22_X1 port map( A1 => n11321, A2 => n11533, B1 => n8644, B2 => 
                           n10529, ZN => n1931);
   U8703 : OAI22_X1 port map( A1 => n11321, A2 => n11541, B1 => n8642, B2 => 
                           n10529, ZN => n1933);
   U8704 : OAI22_X1 port map( A1 => n11321, A2 => n11545, B1 => n8641, B2 => 
                           n11436, ZN => n1934);
   U8705 : OAI22_X1 port map( A1 => n11321, A2 => n11549, B1 => n8640, B2 => 
                           n11436, ZN => n1935);
   U8706 : OAI22_X1 port map( A1 => n11321, A2 => n11553, B1 => n8639, B2 => 
                           n11436, ZN => n1936);
   U8707 : OAI22_X1 port map( A1 => n11321, A2 => n11557, B1 => n8638, B2 => 
                           n11436, ZN => n1937);
   U8708 : OAI22_X1 port map( A1 => n11320, A2 => n11561, B1 => n8637, B2 => 
                           n11436, ZN => n1938);
   U8709 : OAI22_X1 port map( A1 => n11325, A2 => n11493, B1 => n8622, B2 => 
                           n11440, ZN => n1953);
   U8710 : OAI22_X1 port map( A1 => n11325, A2 => n11497, B1 => n8621, B2 => 
                           n11440, ZN => n1954);
   U8711 : OAI22_X1 port map( A1 => n11325, A2 => n11501, B1 => n8620, B2 => 
                           n11440, ZN => n1955);
   U8712 : OAI22_X1 port map( A1 => n11325, A2 => n11505, B1 => n8619, B2 => 
                           n11440, ZN => n1956);
   U8713 : OAI22_X1 port map( A1 => n11325, A2 => n11509, B1 => n8618, B2 => 
                           n11440, ZN => n1957);
   U8714 : OAI22_X1 port map( A1 => n11324, A2 => n11513, B1 => n8617, B2 => 
                           n11440, ZN => n1958);
   U8715 : OAI22_X1 port map( A1 => n11324, A2 => n11517, B1 => n8616, B2 => 
                           n11440, ZN => n1959);
   U8716 : OAI22_X1 port map( A1 => n11324, A2 => n11521, B1 => n8615, B2 => 
                           n11440, ZN => n1960);
   U8717 : OAI22_X1 port map( A1 => n11324, A2 => n11525, B1 => n8614, B2 => 
                           n11440, ZN => n1961);
   U8718 : OAI22_X1 port map( A1 => n11324, A2 => n11529, B1 => n8613, B2 => 
                           n10528, ZN => n1962);
   U8719 : OAI22_X1 port map( A1 => n11324, A2 => n11533, B1 => n8612, B2 => 
                           n10528, ZN => n1963);
   U8720 : OAI22_X1 port map( A1 => n11324, A2 => n11541, B1 => n8610, B2 => 
                           n10528, ZN => n1965);
   U8721 : OAI22_X1 port map( A1 => n11324, A2 => n11545, B1 => n8609, B2 => 
                           n11440, ZN => n1966);
   U8722 : OAI22_X1 port map( A1 => n11324, A2 => n11549, B1 => n8608, B2 => 
                           n11440, ZN => n1967);
   U8723 : OAI22_X1 port map( A1 => n11324, A2 => n11553, B1 => n8607, B2 => 
                           n11440, ZN => n1968);
   U8724 : OAI22_X1 port map( A1 => n11324, A2 => n11557, B1 => n8606, B2 => 
                           n11440, ZN => n1969);
   U8725 : OAI22_X1 port map( A1 => n11323, A2 => n11561, B1 => n8605, B2 => 
                           n11440, ZN => n1970);
   U8726 : OAI22_X1 port map( A1 => n11323, A2 => n11565, B1 => n8604, B2 => 
                           n11440, ZN => n1971);
   U8727 : OAI22_X1 port map( A1 => n11323, A2 => n11569, B1 => n8603, B2 => 
                           n11440, ZN => n1972);
   U8728 : OAI22_X1 port map( A1 => n11323, A2 => n11573, B1 => n8602, B2 => 
                           n11440, ZN => n1973);
   U8729 : OAI22_X1 port map( A1 => n11323, A2 => n11577, B1 => n8601, B2 => 
                           n10528, ZN => n1974);
   U8730 : OAI22_X1 port map( A1 => n11323, A2 => n11581, B1 => n8600, B2 => 
                           n10528, ZN => n1975);
   U8731 : OAI22_X1 port map( A1 => n11323, A2 => n11585, B1 => n8599, B2 => 
                           n10528, ZN => n1976);
   U8732 : OAI22_X1 port map( A1 => n11323, A2 => n11589, B1 => n8598, B2 => 
                           n10528, ZN => n1977);
   U8733 : OAI22_X1 port map( A1 => n11323, A2 => n11593, B1 => n8597, B2 => 
                           n10528, ZN => n1978);
   U8734 : OAI22_X1 port map( A1 => n11323, A2 => n11597, B1 => n8596, B2 => 
                           n10528, ZN => n1979);
   U8735 : OAI22_X1 port map( A1 => n11323, A2 => n11601, B1 => n8595, B2 => 
                           n10528, ZN => n1980);
   U8736 : OAI22_X1 port map( A1 => n11323, A2 => n11609, B1 => n8594, B2 => 
                           n10528, ZN => n1981);
   U8737 : OAI22_X1 port map( A1 => n11340, A2 => n11481, B1 => n8465, B2 => 
                           n11460, ZN => n2110);
   U8738 : OAI22_X1 port map( A1 => n11340, A2 => n11485, B1 => n8464, B2 => 
                           n11460, ZN => n2111);
   U8739 : OAI22_X1 port map( A1 => n11340, A2 => n11489, B1 => n8463, B2 => 
                           n11460, ZN => n2112);
   U8740 : OAI22_X1 port map( A1 => n11340, A2 => n11493, B1 => n8462, B2 => 
                           n11460, ZN => n2113);
   U8741 : OAI22_X1 port map( A1 => n11340, A2 => n11497, B1 => n8461, B2 => 
                           n11460, ZN => n2114);
   U8742 : OAI22_X1 port map( A1 => n11340, A2 => n11501, B1 => n8460, B2 => 
                           n11460, ZN => n2115);
   U8743 : OAI22_X1 port map( A1 => n11340, A2 => n11505, B1 => n8459, B2 => 
                           n11460, ZN => n2116);
   U8744 : OAI22_X1 port map( A1 => n11340, A2 => n11509, B1 => n8458, B2 => 
                           n11460, ZN => n2117);
   U8745 : OAI22_X1 port map( A1 => n11339, A2 => n11513, B1 => n8457, B2 => 
                           n11460, ZN => n2118);
   U8746 : OAI22_X1 port map( A1 => n11339, A2 => n11517, B1 => n8456, B2 => 
                           n11460, ZN => n2119);
   U8747 : OAI22_X1 port map( A1 => n11339, A2 => n11521, B1 => n8455, B2 => 
                           n11460, ZN => n2120);
   U8748 : OAI22_X1 port map( A1 => n11339, A2 => n11557, B1 => n8446, B2 => 
                           n10522, ZN => n2129);
   U8749 : OAI22_X1 port map( A1 => n11338, A2 => n11561, B1 => n8445, B2 => 
                           n10522, ZN => n2130);
   U8750 : OAI22_X1 port map( A1 => n11338, A2 => n11565, B1 => n8444, B2 => 
                           n10522, ZN => n2131);
   U8751 : OAI22_X1 port map( A1 => n11338, A2 => n11569, B1 => n8443, B2 => 
                           n11460, ZN => n2132);
   U8752 : OAI22_X1 port map( A1 => n11338, A2 => n11573, B1 => n8442, B2 => 
                           n11460, ZN => n2133);
   U8753 : OAI22_X1 port map( A1 => n11338, A2 => n11577, B1 => n8441, B2 => 
                           n10522, ZN => n2134);
   U8754 : OAI22_X1 port map( A1 => n11338, A2 => n11581, B1 => n8440, B2 => 
                           n10522, ZN => n2135);
   U8755 : OAI22_X1 port map( A1 => n11338, A2 => n11585, B1 => n8439, B2 => 
                           n10522, ZN => n2136);
   U8756 : OAI22_X1 port map( A1 => n11338, A2 => n11589, B1 => n8438, B2 => 
                           n10522, ZN => n2137);
   U8757 : OAI22_X1 port map( A1 => n11338, A2 => n11593, B1 => n8437, B2 => 
                           n10522, ZN => n2138);
   U8758 : OAI22_X1 port map( A1 => n11338, A2 => n11597, B1 => n8436, B2 => 
                           n10522, ZN => n2139);
   U8759 : OAI22_X1 port map( A1 => n11338, A2 => n11601, B1 => n8435, B2 => 
                           n10522, ZN => n2140);
   U8760 : OAI22_X1 port map( A1 => n11338, A2 => n11609, B1 => n8434, B2 => 
                           n10522, ZN => n2141);
   U8761 : OAI22_X1 port map( A1 => n11348, A2 => n11513, B1 => n8361, B2 => 
                           n11472, ZN => n2214);
   U8762 : OAI22_X1 port map( A1 => n11348, A2 => n11557, B1 => n8350, B2 => 
                           n11472, ZN => n2225);
   U8763 : OAI22_X1 port map( A1 => n11347, A2 => n11565, B1 => n8348, B2 => 
                           n11472, ZN => n2227);
   U8764 : OAI22_X1 port map( A1 => n11347, A2 => n11569, B1 => n8347, B2 => 
                           n11472, ZN => n2228);
   U8765 : OAI22_X1 port map( A1 => n11347, A2 => n11577, B1 => n8345, B2 => 
                           n10515, ZN => n2230);
   U8766 : OAI22_X1 port map( A1 => n11347, A2 => n11585, B1 => n8343, B2 => 
                           n10515, ZN => n2232);
   U8767 : OAI22_X1 port map( A1 => n11322, A2 => n11489, B1 => n8655, B2 => 
                           n11436, ZN => n1920);
   U8768 : OAI22_X1 port map( A1 => n11321, A2 => n11537, B1 => n8643, B2 => 
                           n11436, ZN => n1932);
   U8769 : OAI22_X1 port map( A1 => n11320, A2 => n11565, B1 => n8636, B2 => 
                           n11436, ZN => n1939);
   U8770 : OAI22_X1 port map( A1 => n11320, A2 => n11569, B1 => n8635, B2 => 
                           n11436, ZN => n1940);
   U8771 : OAI22_X1 port map( A1 => n11320, A2 => n11573, B1 => n8634, B2 => 
                           n11436, ZN => n1941);
   U8772 : OAI22_X1 port map( A1 => n11320, A2 => n11577, B1 => n8633, B2 => 
                           n10529, ZN => n1942);
   U8773 : OAI22_X1 port map( A1 => n11320, A2 => n11581, B1 => n8632, B2 => 
                           n10529, ZN => n1943);
   U8774 : OAI22_X1 port map( A1 => n11320, A2 => n11585, B1 => n8631, B2 => 
                           n10529, ZN => n1944);
   U8775 : OAI22_X1 port map( A1 => n11320, A2 => n11589, B1 => n8630, B2 => 
                           n10529, ZN => n1945);
   U8776 : OAI22_X1 port map( A1 => n11320, A2 => n11593, B1 => n8629, B2 => 
                           n10529, ZN => n1946);
   U8777 : OAI22_X1 port map( A1 => n11320, A2 => n11597, B1 => n8628, B2 => 
                           n10529, ZN => n1947);
   U8778 : OAI22_X1 port map( A1 => n11320, A2 => n11601, B1 => n8627, B2 => 
                           n10529, ZN => n1948);
   U8779 : OAI22_X1 port map( A1 => n11320, A2 => n11609, B1 => n8626, B2 => 
                           n10529, ZN => n1949);
   U8780 : OAI22_X1 port map( A1 => n11325, A2 => n11481, B1 => n8625, B2 => 
                           n11440, ZN => n1950);
   U8781 : OAI22_X1 port map( A1 => n11325, A2 => n11485, B1 => n8624, B2 => 
                           n11440, ZN => n1951);
   U8782 : OAI22_X1 port map( A1 => n11325, A2 => n11489, B1 => n8623, B2 => 
                           n11440, ZN => n1952);
   U8783 : OAI22_X1 port map( A1 => n11324, A2 => n11537, B1 => n8611, B2 => 
                           n11440, ZN => n1964);
   U8784 : OAI22_X1 port map( A1 => n11339, A2 => n11525, B1 => n8454, B2 => 
                           n11460, ZN => n2121);
   U8785 : OAI22_X1 port map( A1 => n11339, A2 => n11529, B1 => n8453, B2 => 
                           n11460, ZN => n2122);
   U8786 : OAI22_X1 port map( A1 => n11339, A2 => n11533, B1 => n8452, B2 => 
                           n11460, ZN => n2123);
   U8787 : OAI22_X1 port map( A1 => n11339, A2 => n11537, B1 => n8451, B2 => 
                           n11460, ZN => n2124);
   U8788 : OAI22_X1 port map( A1 => n11339, A2 => n11541, B1 => n8450, B2 => 
                           n11460, ZN => n2125);
   U8789 : OAI22_X1 port map( A1 => n11339, A2 => n11545, B1 => n8449, B2 => 
                           n11460, ZN => n2126);
   U8790 : OAI22_X1 port map( A1 => n11339, A2 => n11549, B1 => n8448, B2 => 
                           n11460, ZN => n2127);
   U8791 : OAI22_X1 port map( A1 => n11339, A2 => n11553, B1 => n8447, B2 => 
                           n11460, ZN => n2128);
   U8792 : OAI22_X1 port map( A1 => n11352, A2 => n11481, B1 => n8337, B2 => 
                           n11476, ZN => n2238);
   U8793 : OAI22_X1 port map( A1 => n11352, A2 => n11485, B1 => n8336, B2 => 
                           n11476, ZN => n2239);
   U8794 : OAI22_X1 port map( A1 => n11352, A2 => n11489, B1 => n8335, B2 => 
                           n11476, ZN => n2240);
   U8795 : OAI22_X1 port map( A1 => n11352, A2 => n11493, B1 => n8334, B2 => 
                           n11476, ZN => n2241);
   U8796 : OAI22_X1 port map( A1 => n11352, A2 => n11497, B1 => n8333, B2 => 
                           n11476, ZN => n2242);
   U8797 : OAI22_X1 port map( A1 => n11352, A2 => n11501, B1 => n8332, B2 => 
                           n11476, ZN => n2243);
   U8798 : OAI22_X1 port map( A1 => n11352, A2 => n11505, B1 => n8331, B2 => 
                           n11476, ZN => n2244);
   U8799 : OAI22_X1 port map( A1 => n11352, A2 => n11509, B1 => n8330, B2 => 
                           n11476, ZN => n2245);
   U8800 : OAI22_X1 port map( A1 => n11351, A2 => n11513, B1 => n8329, B2 => 
                           n11476, ZN => n2246);
   U8801 : OAI22_X1 port map( A1 => n11351, A2 => n11517, B1 => n8328, B2 => 
                           n11476, ZN => n2247);
   U8802 : OAI22_X1 port map( A1 => n11351, A2 => n11521, B1 => n8327, B2 => 
                           n11476, ZN => n2248);
   U8803 : OAI22_X1 port map( A1 => n11351, A2 => n11525, B1 => n8326, B2 => 
                           n11476, ZN => n2249);
   U8804 : OAI22_X1 port map( A1 => n11351, A2 => n11529, B1 => n8325, B2 => 
                           n10513, ZN => n2250);
   U8805 : OAI22_X1 port map( A1 => n11351, A2 => n11533, B1 => n8324, B2 => 
                           n10513, ZN => n2251);
   U8806 : OAI22_X1 port map( A1 => n11351, A2 => n11537, B1 => n8323, B2 => 
                           n10513, ZN => n2252);
   U8807 : OAI22_X1 port map( A1 => n11351, A2 => n11541, B1 => n8322, B2 => 
                           n11476, ZN => n2253);
   U8808 : OAI22_X1 port map( A1 => n11351, A2 => n11545, B1 => n8321, B2 => 
                           n11476, ZN => n2254);
   U8809 : OAI22_X1 port map( A1 => n11351, A2 => n11549, B1 => n8320, B2 => 
                           n11476, ZN => n2255);
   U8810 : OAI22_X1 port map( A1 => n11351, A2 => n11553, B1 => n8319, B2 => 
                           n11476, ZN => n2256);
   U8811 : OAI22_X1 port map( A1 => n11351, A2 => n11557, B1 => n8318, B2 => 
                           n11476, ZN => n2257);
   U8812 : OAI22_X1 port map( A1 => n11350, A2 => n11561, B1 => n8317, B2 => 
                           n11476, ZN => n2258);
   U8813 : OAI22_X1 port map( A1 => n11350, A2 => n11565, B1 => n8316, B2 => 
                           n11476, ZN => n2259);
   U8814 : OAI22_X1 port map( A1 => n11350, A2 => n11569, B1 => n8315, B2 => 
                           n11476, ZN => n2260);
   U8815 : OAI22_X1 port map( A1 => n11350, A2 => n11573, B1 => n8314, B2 => 
                           n11476, ZN => n2261);
   U8816 : OAI22_X1 port map( A1 => n11350, A2 => n11577, B1 => n8313, B2 => 
                           n10513, ZN => n2262);
   U8817 : OAI22_X1 port map( A1 => n11350, A2 => n11581, B1 => n8312, B2 => 
                           n10513, ZN => n2263);
   U8818 : OAI22_X1 port map( A1 => n11350, A2 => n11585, B1 => n8311, B2 => 
                           n10513, ZN => n2264);
   U8819 : OAI22_X1 port map( A1 => n11350, A2 => n11589, B1 => n8310, B2 => 
                           n10513, ZN => n2265);
   U8820 : OAI22_X1 port map( A1 => n11350, A2 => n11593, B1 => n8309, B2 => 
                           n10513, ZN => n2266);
   U8821 : OAI22_X1 port map( A1 => n11350, A2 => n11597, B1 => n8308, B2 => 
                           n10513, ZN => n2267);
   U8822 : OAI22_X1 port map( A1 => n11350, A2 => n11601, B1 => n8307, B2 => 
                           n10513, ZN => n2268);
   U8823 : OAI22_X1 port map( A1 => n11350, A2 => n11609, B1 => n8306, B2 => 
                           n10513, ZN => n2269);
   U8824 : OAI22_X1 port map( A1 => n9297, A2 => n11356, B1 => n11262, B2 => 
                           n11483, ZN => n1278);
   U8825 : OAI22_X1 port map( A1 => n9296, A2 => n11356, B1 => n11262, B2 => 
                           n11487, ZN => n1279);
   U8826 : OAI22_X1 port map( A1 => n9295, A2 => n11356, B1 => n11262, B2 => 
                           n11491, ZN => n1280);
   U8827 : OAI22_X1 port map( A1 => n9294, A2 => n11356, B1 => n11262, B2 => 
                           n11495, ZN => n1281);
   U8828 : OAI22_X1 port map( A1 => n9293, A2 => n11356, B1 => n11262, B2 => 
                           n11499, ZN => n1282);
   U8829 : OAI22_X1 port map( A1 => n9292, A2 => n11356, B1 => n11262, B2 => 
                           n11503, ZN => n1283);
   U8830 : OAI22_X1 port map( A1 => n9291, A2 => n11356, B1 => n11262, B2 => 
                           n11507, ZN => n1284);
   U8831 : OAI22_X1 port map( A1 => n9290, A2 => n11356, B1 => n11262, B2 => 
                           n11511, ZN => n1285);
   U8832 : OAI22_X1 port map( A1 => n9289, A2 => n11356, B1 => n11261, B2 => 
                           n11515, ZN => n1286);
   U8833 : OAI22_X1 port map( A1 => n9288, A2 => n11356, B1 => n11261, B2 => 
                           n11519, ZN => n1287);
   U8834 : OAI22_X1 port map( A1 => n9287, A2 => n11356, B1 => n11261, B2 => 
                           n11523, ZN => n1288);
   U8835 : OAI22_X1 port map( A1 => n9286, A2 => n11356, B1 => n11261, B2 => 
                           n11527, ZN => n1289);
   U8836 : OAI22_X1 port map( A1 => n9285, A2 => n10555, B1 => n11261, B2 => 
                           n11531, ZN => n1290);
   U8837 : OAI22_X1 port map( A1 => n9284, A2 => n10555, B1 => n11261, B2 => 
                           n11535, ZN => n1291);
   U8838 : OAI22_X1 port map( A1 => n9283, A2 => n10555, B1 => n11261, B2 => 
                           n11539, ZN => n1292);
   U8839 : OAI22_X1 port map( A1 => n9282, A2 => n11356, B1 => n11261, B2 => 
                           n11543, ZN => n1293);
   U8840 : OAI22_X1 port map( A1 => n9281, A2 => n11356, B1 => n11261, B2 => 
                           n11547, ZN => n1294);
   U8841 : OAI22_X1 port map( A1 => n9280, A2 => n11356, B1 => n11261, B2 => 
                           n11551, ZN => n1295);
   U8842 : OAI22_X1 port map( A1 => n9279, A2 => n11356, B1 => n11261, B2 => 
                           n11555, ZN => n1296);
   U8843 : OAI22_X1 port map( A1 => n9278, A2 => n11356, B1 => n11261, B2 => 
                           n11559, ZN => n1297);
   U8844 : OAI22_X1 port map( A1 => n9277, A2 => n11356, B1 => n11260, B2 => 
                           n11563, ZN => n1298);
   U8845 : OAI22_X1 port map( A1 => n9276, A2 => n11356, B1 => n11260, B2 => 
                           n11567, ZN => n1299);
   U8846 : OAI22_X1 port map( A1 => n9275, A2 => n11356, B1 => n11260, B2 => 
                           n11571, ZN => n1300);
   U8847 : OAI22_X1 port map( A1 => n9274, A2 => n11356, B1 => n11260, B2 => 
                           n11575, ZN => n1301);
   U8848 : OAI22_X1 port map( A1 => n9273, A2 => n10555, B1 => n11260, B2 => 
                           n11579, ZN => n1302);
   U8849 : OAI22_X1 port map( A1 => n9272, A2 => n10555, B1 => n11260, B2 => 
                           n11583, ZN => n1303);
   U8850 : OAI22_X1 port map( A1 => n9271, A2 => n10555, B1 => n11260, B2 => 
                           n11587, ZN => n1304);
   U8851 : OAI22_X1 port map( A1 => n9270, A2 => n10555, B1 => n11260, B2 => 
                           n11591, ZN => n1305);
   U8852 : OAI22_X1 port map( A1 => n9269, A2 => n10555, B1 => n11260, B2 => 
                           n11595, ZN => n1306);
   U8853 : OAI22_X1 port map( A1 => n9268, A2 => n10555, B1 => n11260, B2 => 
                           n11599, ZN => n1307);
   U8854 : OAI22_X1 port map( A1 => n9267, A2 => n10555, B1 => n11260, B2 => 
                           n11603, ZN => n1308);
   U8855 : OAI22_X1 port map( A1 => n9266, A2 => n10555, B1 => n11260, B2 => 
                           n11611, ZN => n1309);
   U8856 : NOR3_X1 port map( A1 => n8272, A2 => n8273, A3 => n8271, ZN => 
                           n10458);
   U8857 : NOR3_X1 port map( A1 => n8268, A2 => n8269, A3 => n8267, ZN => n9868
                           );
   U8858 : NAND2_X1 port map( A1 => n8264, A2 => n8265, ZN => n10512);
   U8859 : NAND2_X1 port map( A1 => n10472, A2 => n10454, ZN => n9922);
   U8860 : NAND2_X1 port map( A1 => n10473, A2 => n10472, ZN => n9921);
   U8861 : NAND2_X1 port map( A1 => n10474, A2 => n10473, ZN => n9920);
   U8862 : NAND2_X1 port map( A1 => n10474, A2 => n10463, ZN => n9933);
   U8863 : NAND2_X1 port map( A1 => n10474, A2 => n10460, ZN => n9932);
   U8864 : NAND2_X1 port map( A1 => n10472, A2 => n10463, ZN => n9931);
   U8865 : NAND2_X1 port map( A1 => n10472, A2 => n10460, ZN => n9926);
   U8866 : NAND2_X1 port map( A1 => n10474, A2 => n10456, ZN => n9927);
   U8867 : NAND2_X1 port map( A1 => n10473, A2 => n10455, ZN => n9937);
   U8868 : NAND2_X1 port map( A1 => n10473, A2 => n10457, ZN => n9938);
   U8869 : NAND2_X1 port map( A1 => n9882, A2 => n9864, ZN => n9332);
   U8870 : NAND2_X1 port map( A1 => n9883, A2 => n9882, ZN => n9331);
   U8871 : NAND2_X1 port map( A1 => n9884, A2 => n9883, ZN => n9330);
   U8872 : NAND2_X1 port map( A1 => n9884, A2 => n9873, ZN => n9343);
   U8873 : NAND2_X1 port map( A1 => n9884, A2 => n9870, ZN => n9342);
   U8874 : NAND2_X1 port map( A1 => n9882, A2 => n9873, ZN => n9341);
   U8875 : NAND2_X1 port map( A1 => n9884, A2 => n9866, ZN => n9337);
   U8876 : NAND2_X1 port map( A1 => n9882, A2 => n9870, ZN => n9336);
   U8877 : NAND2_X1 port map( A1 => n9883, A2 => n9867, ZN => n9348);
   U8878 : NAND2_X1 port map( A1 => n9883, A2 => n9865, ZN => n9347);
   U8879 : AND3_X1 port map( A1 => n10454, A2 => n11698, A3 => n10457, ZN => 
                           n9892);
   U8880 : AND3_X1 port map( A1 => n10455, A2 => n11698, A3 => n10463, ZN => 
                           n9902);
   U8881 : AND3_X1 port map( A1 => n9864, A2 => n11837, A3 => n9867, ZN => 
                           n9302);
   U8882 : AND3_X1 port map( A1 => n9865, A2 => n11837, A3 => n9873, ZN => 
                           n9312);
   U8883 : AND3_X1 port map( A1 => n10457, A2 => n11698, A3 => n10458, ZN => 
                           n9893);
   U8884 : AND3_X1 port map( A1 => n10457, A2 => n11698, A3 => n10461, ZN => 
                           n9897);
   U8885 : AND3_X1 port map( A1 => n10455, A2 => n11698, A3 => n10456, ZN => 
                           n9898);
   U8886 : AND3_X1 port map( A1 => n10455, A2 => n11698, A3 => n10464, ZN => 
                           n9903);
   U8887 : AND3_X1 port map( A1 => n9867, A2 => n11837, A3 => n9868, ZN => 
                           n9303);
   U8888 : AND3_X1 port map( A1 => n9865, A2 => n11837, A3 => n9866, ZN => 
                           n9308);
   U8889 : AND3_X1 port map( A1 => n9867, A2 => n11837, A3 => n9871, ZN => 
                           n9307);
   U8890 : AND3_X1 port map( A1 => n9865, A2 => n11837, A3 => n9874, ZN => 
                           n9313);
   U8891 : AND2_X1 port map( A1 => n10474, A2 => n10454, ZN => n9917);
   U8892 : AND2_X1 port map( A1 => n10472, A2 => n10458, ZN => n9918);
   U8893 : AND2_X1 port map( A1 => n10472, A2 => n10461, ZN => n9928);
   U8894 : AND2_X1 port map( A1 => n10474, A2 => n10461, ZN => n9929);
   U8895 : AND2_X1 port map( A1 => n10474, A2 => n10458, ZN => n9923);
   U8896 : AND2_X1 port map( A1 => n10472, A2 => n10456, ZN => n9924);
   U8897 : AND2_X1 port map( A1 => n10472, A2 => n10464, ZN => n9934);
   U8898 : AND2_X1 port map( A1 => n10474, A2 => n10464, ZN => n9935);
   U8899 : AND2_X1 port map( A1 => n9882, A2 => n9868, ZN => n9328);
   U8900 : AND2_X1 port map( A1 => n9884, A2 => n9864, ZN => n9327);
   U8901 : AND2_X1 port map( A1 => n9884, A2 => n9871, ZN => n9339);
   U8902 : AND2_X1 port map( A1 => n9882, A2 => n9871, ZN => n9338);
   U8903 : AND2_X1 port map( A1 => n9882, A2 => n9866, ZN => n9334);
   U8904 : AND2_X1 port map( A1 => n9884, A2 => n9868, ZN => n9333);
   U8905 : AND2_X1 port map( A1 => n9884, A2 => n9874, ZN => n9345);
   U8906 : AND2_X1 port map( A1 => n9882, A2 => n9874, ZN => n9344);
   U8907 : INV_X1 port map( A => n10555, ZN => n11359);
   U8908 : OAI21_X1 port map( B1 => n10518, B2 => n10552, A => n11895, ZN => 
                           n10555);
   U8909 : INV_X1 port map( A => n10554, ZN => n11363);
   U8910 : OAI21_X1 port map( B1 => n10516, B2 => n10552, A => n11892, ZN => 
                           n10554);
   U8911 : INV_X1 port map( A => n10553, ZN => n11367);
   U8912 : OAI21_X1 port map( B1 => n10514, B2 => n10552, A => n11892, ZN => 
                           n10553);
   U8913 : INV_X1 port map( A => n10551, ZN => n11371);
   U8914 : OAI21_X1 port map( B1 => n10512, B2 => n10552, A => n11892, ZN => 
                           n10551);
   U8915 : INV_X1 port map( A => n10550, ZN => n11375);
   U8916 : OAI21_X1 port map( B1 => n10518, B2 => n10547, A => n11893, ZN => 
                           n10550);
   U8917 : INV_X1 port map( A => n10549, ZN => n11379);
   U8918 : OAI21_X1 port map( B1 => n10516, B2 => n10547, A => n11893, ZN => 
                           n10549);
   U8919 : INV_X1 port map( A => n10548, ZN => n11383);
   U8920 : OAI21_X1 port map( B1 => n10514, B2 => n10547, A => n11893, ZN => 
                           n10548);
   U8921 : INV_X1 port map( A => n10546, ZN => n11387);
   U8922 : OAI21_X1 port map( B1 => n10512, B2 => n10547, A => n11893, ZN => 
                           n10546);
   U8923 : INV_X1 port map( A => n10545, ZN => n11391);
   U8924 : OAI21_X1 port map( B1 => n10518, B2 => n10542, A => n11893, ZN => 
                           n10545);
   U8925 : INV_X1 port map( A => n10544, ZN => n11395);
   U8926 : OAI21_X1 port map( B1 => n10516, B2 => n10542, A => n11893, ZN => 
                           n10544);
   U8927 : INV_X1 port map( A => n10543, ZN => n11399);
   U8928 : OAI21_X1 port map( B1 => n10514, B2 => n10542, A => n11893, ZN => 
                           n10543);
   U8929 : INV_X1 port map( A => n10541, ZN => n11403);
   U8930 : OAI21_X1 port map( B1 => n10512, B2 => n10542, A => n11893, ZN => 
                           n10541);
   U8931 : INV_X1 port map( A => n10539, ZN => n11407);
   U8932 : OAI21_X1 port map( B1 => n10518, B2 => n10536, A => n11893, ZN => 
                           n10539);
   U8933 : INV_X1 port map( A => n10538, ZN => n11411);
   U8934 : OAI21_X1 port map( B1 => n10516, B2 => n10536, A => n11893, ZN => 
                           n10538);
   U8935 : INV_X1 port map( A => n10537, ZN => n11415);
   U8936 : OAI21_X1 port map( B1 => n10514, B2 => n10536, A => n11893, ZN => 
                           n10537);
   U8937 : INV_X1 port map( A => n10534, ZN => n11423);
   U8938 : OAI21_X1 port map( B1 => n10518, B2 => n10531, A => n11893, ZN => 
                           n10534);
   U8939 : INV_X1 port map( A => n10533, ZN => n11427);
   U8940 : OAI21_X1 port map( B1 => n10516, B2 => n10531, A => n11894, ZN => 
                           n10533);
   U8941 : INV_X1 port map( A => n10532, ZN => n11431);
   U8942 : OAI21_X1 port map( B1 => n10514, B2 => n10531, A => n11894, ZN => 
                           n10532);
   U8943 : INV_X1 port map( A => n10530, ZN => n11435);
   U8944 : OAI21_X1 port map( B1 => n10512, B2 => n10531, A => n11894, ZN => 
                           n10530);
   U8945 : INV_X1 port map( A => n10529, ZN => n11439);
   U8946 : OAI21_X1 port map( B1 => n10518, B2 => n10526, A => n11894, ZN => 
                           n10529);
   U8947 : INV_X1 port map( A => n10528, ZN => n11443);
   U8948 : OAI21_X1 port map( B1 => n10516, B2 => n10526, A => n11894, ZN => 
                           n10528);
   U8949 : INV_X1 port map( A => n10527, ZN => n11447);
   U8950 : OAI21_X1 port map( B1 => n10514, B2 => n10526, A => n11894, ZN => 
                           n10527);
   U8951 : INV_X1 port map( A => n10525, ZN => n11451);
   U8952 : OAI21_X1 port map( B1 => n10512, B2 => n10526, A => n11894, ZN => 
                           n10525);
   U8953 : INV_X1 port map( A => n10524, ZN => n11455);
   U8954 : OAI21_X1 port map( B1 => n10518, B2 => n10521, A => n11894, ZN => 
                           n10524);
   U8955 : INV_X1 port map( A => n10523, ZN => n11459);
   U8956 : OAI21_X1 port map( B1 => n10516, B2 => n10521, A => n11894, ZN => 
                           n10523);
   U8957 : INV_X1 port map( A => n10522, ZN => n11463);
   U8958 : OAI21_X1 port map( B1 => n10514, B2 => n10521, A => n11894, ZN => 
                           n10522);
   U8959 : INV_X1 port map( A => n10520, ZN => n11467);
   U8960 : OAI21_X1 port map( B1 => n10512, B2 => n10521, A => n11894, ZN => 
                           n10520);
   U8961 : INV_X1 port map( A => n10517, ZN => n11471);
   U8962 : OAI21_X1 port map( B1 => n10511, B2 => n10518, A => n11894, ZN => 
                           n10517);
   U8963 : INV_X1 port map( A => n10515, ZN => n11475);
   U8964 : OAI21_X1 port map( B1 => n10511, B2 => n10516, A => n11894, ZN => 
                           n10515);
   U8965 : INV_X1 port map( A => n10513, ZN => n11479);
   U8966 : OAI21_X1 port map( B1 => n10511, B2 => n10514, A => n11895, ZN => 
                           n10513);
   U8967 : BUF_X1 port map( A => n11695, Z => n11692);
   U8968 : BUF_X1 port map( A => n11834, Z => n11831);
   U8969 : BUF_X1 port map( A => n11695, Z => n11693);
   U8970 : BUF_X1 port map( A => n11834, Z => n11832);
   U8971 : BUF_X1 port map( A => n11480, Z => n11482);
   U8972 : BUF_X1 port map( A => n11484, Z => n11486);
   U8973 : BUF_X1 port map( A => n11488, Z => n11490);
   U8974 : BUF_X1 port map( A => n11492, Z => n11494);
   U8975 : BUF_X1 port map( A => n11496, Z => n11498);
   U8976 : BUF_X1 port map( A => n11500, Z => n11502);
   U8977 : BUF_X1 port map( A => n11504, Z => n11506);
   U8978 : BUF_X1 port map( A => n11508, Z => n11510);
   U8979 : BUF_X1 port map( A => n11512, Z => n11514);
   U8980 : BUF_X1 port map( A => n11516, Z => n11518);
   U8981 : BUF_X1 port map( A => n11520, Z => n11522);
   U8982 : BUF_X1 port map( A => n11524, Z => n11526);
   U8983 : BUF_X1 port map( A => n11528, Z => n11530);
   U8984 : BUF_X1 port map( A => n11532, Z => n11534);
   U8985 : BUF_X1 port map( A => n11536, Z => n11538);
   U8986 : BUF_X1 port map( A => n11540, Z => n11542);
   U8987 : BUF_X1 port map( A => n11544, Z => n11546);
   U8988 : BUF_X1 port map( A => n11548, Z => n11550);
   U8989 : BUF_X1 port map( A => n11552, Z => n11554);
   U8990 : BUF_X1 port map( A => n11556, Z => n11558);
   U8991 : BUF_X1 port map( A => n11560, Z => n11562);
   U8992 : BUF_X1 port map( A => n11564, Z => n11566);
   U8993 : BUF_X1 port map( A => n11568, Z => n11570);
   U8994 : BUF_X1 port map( A => n11572, Z => n11574);
   U8995 : BUF_X1 port map( A => n11576, Z => n11578);
   U8996 : BUF_X1 port map( A => n11580, Z => n11582);
   U8997 : BUF_X1 port map( A => n11584, Z => n11586);
   U8998 : BUF_X1 port map( A => n11588, Z => n11590);
   U8999 : BUF_X1 port map( A => n11592, Z => n11594);
   U9000 : BUF_X1 port map( A => n11596, Z => n11598);
   U9001 : BUF_X1 port map( A => n11600, Z => n11602);
   U9002 : BUF_X1 port map( A => n11608, Z => n11610);
   U9003 : BUF_X1 port map( A => n11480, Z => n11481);
   U9004 : BUF_X1 port map( A => n11484, Z => n11485);
   U9005 : BUF_X1 port map( A => n11488, Z => n11489);
   U9006 : BUF_X1 port map( A => n11492, Z => n11493);
   U9007 : BUF_X1 port map( A => n11496, Z => n11497);
   U9008 : BUF_X1 port map( A => n11500, Z => n11501);
   U9009 : BUF_X1 port map( A => n11504, Z => n11505);
   U9010 : BUF_X1 port map( A => n11508, Z => n11509);
   U9011 : BUF_X1 port map( A => n11512, Z => n11513);
   U9012 : BUF_X1 port map( A => n11516, Z => n11517);
   U9013 : BUF_X1 port map( A => n11520, Z => n11521);
   U9014 : BUF_X1 port map( A => n11524, Z => n11525);
   U9015 : BUF_X1 port map( A => n11528, Z => n11529);
   U9016 : BUF_X1 port map( A => n11532, Z => n11533);
   U9017 : BUF_X1 port map( A => n11536, Z => n11537);
   U9018 : BUF_X1 port map( A => n11540, Z => n11541);
   U9019 : BUF_X1 port map( A => n11544, Z => n11545);
   U9020 : BUF_X1 port map( A => n11548, Z => n11549);
   U9021 : BUF_X1 port map( A => n11552, Z => n11553);
   U9022 : BUF_X1 port map( A => n11556, Z => n11557);
   U9023 : BUF_X1 port map( A => n11560, Z => n11561);
   U9024 : BUF_X1 port map( A => n11564, Z => n11565);
   U9025 : BUF_X1 port map( A => n11568, Z => n11569);
   U9026 : BUF_X1 port map( A => n11572, Z => n11573);
   U9027 : BUF_X1 port map( A => n11576, Z => n11577);
   U9028 : BUF_X1 port map( A => n11580, Z => n11581);
   U9029 : BUF_X1 port map( A => n11584, Z => n11585);
   U9030 : BUF_X1 port map( A => n11588, Z => n11589);
   U9031 : BUF_X1 port map( A => n11592, Z => n11593);
   U9032 : BUF_X1 port map( A => n11596, Z => n11597);
   U9033 : BUF_X1 port map( A => n11600, Z => n11601);
   U9034 : BUF_X1 port map( A => n11608, Z => n11609);
   U9035 : BUF_X1 port map( A => n11701, Z => n11696);
   U9036 : BUF_X1 port map( A => n11702, Z => n11701);
   U9037 : BUF_X1 port map( A => n11840, Z => n11835);
   U9038 : BUF_X1 port map( A => n11841, Z => n11840);
   U9039 : BUF_X1 port map( A => n11480, Z => n11483);
   U9040 : BUF_X1 port map( A => n11484, Z => n11487);
   U9041 : BUF_X1 port map( A => n11488, Z => n11491);
   U9042 : BUF_X1 port map( A => n11492, Z => n11495);
   U9043 : BUF_X1 port map( A => n11496, Z => n11499);
   U9044 : BUF_X1 port map( A => n11500, Z => n11503);
   U9045 : BUF_X1 port map( A => n11504, Z => n11507);
   U9046 : BUF_X1 port map( A => n11508, Z => n11511);
   U9047 : BUF_X1 port map( A => n11512, Z => n11515);
   U9048 : BUF_X1 port map( A => n11516, Z => n11519);
   U9049 : BUF_X1 port map( A => n11520, Z => n11523);
   U9050 : BUF_X1 port map( A => n11524, Z => n11527);
   U9051 : BUF_X1 port map( A => n11528, Z => n11531);
   U9052 : BUF_X1 port map( A => n11532, Z => n11535);
   U9053 : BUF_X1 port map( A => n11536, Z => n11539);
   U9054 : BUF_X1 port map( A => n11540, Z => n11543);
   U9055 : BUF_X1 port map( A => n11544, Z => n11547);
   U9056 : BUF_X1 port map( A => n11548, Z => n11551);
   U9057 : BUF_X1 port map( A => n11552, Z => n11555);
   U9058 : BUF_X1 port map( A => n11556, Z => n11559);
   U9059 : BUF_X1 port map( A => n11560, Z => n11563);
   U9060 : BUF_X1 port map( A => n11564, Z => n11567);
   U9061 : BUF_X1 port map( A => n11568, Z => n11571);
   U9062 : BUF_X1 port map( A => n11572, Z => n11575);
   U9063 : BUF_X1 port map( A => n11576, Z => n11579);
   U9064 : BUF_X1 port map( A => n11580, Z => n11583);
   U9065 : BUF_X1 port map( A => n11584, Z => n11587);
   U9066 : BUF_X1 port map( A => n11588, Z => n11591);
   U9067 : BUF_X1 port map( A => n11592, Z => n11595);
   U9068 : BUF_X1 port map( A => n11596, Z => n11599);
   U9069 : BUF_X1 port map( A => n11600, Z => n11603);
   U9070 : BUF_X1 port map( A => n11608, Z => n11611);
   U9071 : BUF_X1 port map( A => n11695, Z => n11694);
   U9072 : BUF_X1 port map( A => n11834, Z => n11833);
   U9073 : AOI221_X1 port map( B1 => n10685, B2 => n11820, C1 => n11101, C2 => 
                           n11816, A => n9881, ZN => n9880);
   U9074 : OAI222_X1 port map( A1 => n11812, A2 => n8721, B1 => n11808, B2 => 
                           n8465, C1 => n11804, C2 => n8337, ZN => n9881);
   U9075 : AOI221_X1 port map( B1 => n10686, B2 => n11820, C1 => n11102, C2 => 
                           n11816, A => n9855, ZN => n9854);
   U9076 : OAI222_X1 port map( A1 => n11812, A2 => n8720, B1 => n11808, B2 => 
                           n8464, C1 => n11804, C2 => n8336, ZN => n9855);
   U9077 : AOI221_X1 port map( B1 => n10687, B2 => n11820, C1 => n11103, C2 => 
                           n11816, A => n9838, ZN => n9837);
   U9078 : OAI222_X1 port map( A1 => n11812, A2 => n8719, B1 => n11808, B2 => 
                           n8463, C1 => n11804, C2 => n8335, ZN => n9838);
   U9079 : AOI221_X1 port map( B1 => n10688, B2 => n11820, C1 => n11104, C2 => 
                           n11816, A => n9821, ZN => n9820);
   U9080 : OAI222_X1 port map( A1 => n11812, A2 => n8718, B1 => n11808, B2 => 
                           n8462, C1 => n11804, C2 => n8334, ZN => n9821);
   U9081 : AOI221_X1 port map( B1 => n10689, B2 => n11820, C1 => n11105, C2 => 
                           n11816, A => n9804, ZN => n9803);
   U9082 : OAI222_X1 port map( A1 => n11812, A2 => n8717, B1 => n11808, B2 => 
                           n8461, C1 => n11804, C2 => n8333, ZN => n9804);
   U9083 : AOI221_X1 port map( B1 => n10690, B2 => n11820, C1 => n11106, C2 => 
                           n11816, A => n9787, ZN => n9786);
   U9084 : OAI222_X1 port map( A1 => n11812, A2 => n8716, B1 => n11808, B2 => 
                           n8460, C1 => n11804, C2 => n8332, ZN => n9787);
   U9085 : AOI221_X1 port map( B1 => n10691, B2 => n11820, C1 => n11107, C2 => 
                           n11816, A => n9770, ZN => n9769);
   U9086 : OAI222_X1 port map( A1 => n11812, A2 => n8715, B1 => n11808, B2 => 
                           n8459, C1 => n11804, C2 => n8331, ZN => n9770);
   U9087 : AOI221_X1 port map( B1 => n10692, B2 => n11820, C1 => n11108, C2 => 
                           n11816, A => n9753, ZN => n9752);
   U9088 : OAI222_X1 port map( A1 => n11812, A2 => n8714, B1 => n11808, B2 => 
                           n8458, C1 => n11804, C2 => n8330, ZN => n9753);
   U9089 : AOI221_X1 port map( B1 => n10693, B2 => n11820, C1 => n11109, C2 => 
                           n11816, A => n9736, ZN => n9735);
   U9090 : OAI222_X1 port map( A1 => n11812, A2 => n8713, B1 => n11808, B2 => 
                           n8457, C1 => n11804, C2 => n8329, ZN => n9736);
   U9091 : AOI221_X1 port map( B1 => n10694, B2 => n11820, C1 => n11110, C2 => 
                           n11816, A => n9719, ZN => n9718);
   U9092 : OAI222_X1 port map( A1 => n11812, A2 => n8712, B1 => n11808, B2 => 
                           n8456, C1 => n11804, C2 => n8328, ZN => n9719);
   U9093 : AOI221_X1 port map( B1 => n10695, B2 => n11820, C1 => n11111, C2 => 
                           n11816, A => n9702, ZN => n9701);
   U9094 : OAI222_X1 port map( A1 => n11812, A2 => n8711, B1 => n11808, B2 => 
                           n8455, C1 => n11804, C2 => n8327, ZN => n9702);
   U9095 : AOI221_X1 port map( B1 => n10696, B2 => n11820, C1 => n11112, C2 => 
                           n11816, A => n9685, ZN => n9684);
   U9096 : OAI222_X1 port map( A1 => n11812, A2 => n8710, B1 => n11808, B2 => 
                           n8454, C1 => n11804, C2 => n8326, ZN => n9685);
   U9097 : AOI221_X1 port map( B1 => n10697, B2 => n11821, C1 => n11113, C2 => 
                           n11817, A => n9668, ZN => n9667);
   U9098 : OAI222_X1 port map( A1 => n11813, A2 => n8709, B1 => n11809, B2 => 
                           n8453, C1 => n11805, C2 => n8325, ZN => n9668);
   U9099 : AOI221_X1 port map( B1 => n10698, B2 => n11821, C1 => n11114, C2 => 
                           n11817, A => n9651, ZN => n9650);
   U9100 : OAI222_X1 port map( A1 => n11813, A2 => n8708, B1 => n11809, B2 => 
                           n8452, C1 => n11805, C2 => n8324, ZN => n9651);
   U9101 : AOI221_X1 port map( B1 => n10699, B2 => n11821, C1 => n11115, C2 => 
                           n11817, A => n9634, ZN => n9633);
   U9102 : OAI222_X1 port map( A1 => n11813, A2 => n8707, B1 => n11809, B2 => 
                           n8451, C1 => n11805, C2 => n8323, ZN => n9634);
   U9103 : AOI221_X1 port map( B1 => n10700, B2 => n11821, C1 => n11116, C2 => 
                           n11817, A => n9617, ZN => n9616);
   U9104 : OAI222_X1 port map( A1 => n11813, A2 => n8706, B1 => n11809, B2 => 
                           n8450, C1 => n11805, C2 => n8322, ZN => n9617);
   U9105 : AOI221_X1 port map( B1 => n10701, B2 => n11821, C1 => n11117, C2 => 
                           n11817, A => n9600, ZN => n9599);
   U9106 : OAI222_X1 port map( A1 => n11813, A2 => n8705, B1 => n11809, B2 => 
                           n8449, C1 => n11805, C2 => n8321, ZN => n9600);
   U9107 : AOI221_X1 port map( B1 => n10702, B2 => n11821, C1 => n11118, C2 => 
                           n11817, A => n9583, ZN => n9582);
   U9108 : OAI222_X1 port map( A1 => n11813, A2 => n8704, B1 => n11809, B2 => 
                           n8448, C1 => n11805, C2 => n8320, ZN => n9583);
   U9109 : AOI221_X1 port map( B1 => n10703, B2 => n11821, C1 => n11119, C2 => 
                           n11817, A => n9566, ZN => n9565);
   U9110 : OAI222_X1 port map( A1 => n11813, A2 => n8703, B1 => n11809, B2 => 
                           n8447, C1 => n11805, C2 => n8319, ZN => n9566);
   U9111 : AOI221_X1 port map( B1 => n10704, B2 => n11821, C1 => n11120, C2 => 
                           n11817, A => n9549, ZN => n9548);
   U9112 : OAI222_X1 port map( A1 => n11813, A2 => n8702, B1 => n11809, B2 => 
                           n8446, C1 => n11805, C2 => n8318, ZN => n9549);
   U9113 : AOI221_X1 port map( B1 => n10705, B2 => n11821, C1 => n11121, C2 => 
                           n11817, A => n9532, ZN => n9531);
   U9114 : OAI222_X1 port map( A1 => n11813, A2 => n8701, B1 => n11809, B2 => 
                           n8445, C1 => n11805, C2 => n8317, ZN => n9532);
   U9115 : AOI221_X1 port map( B1 => n10706, B2 => n11821, C1 => n11122, C2 => 
                           n11817, A => n9515, ZN => n9514);
   U9116 : OAI222_X1 port map( A1 => n11813, A2 => n8700, B1 => n11809, B2 => 
                           n8444, C1 => n11805, C2 => n8316, ZN => n9515);
   U9117 : AOI221_X1 port map( B1 => n10707, B2 => n11821, C1 => n11123, C2 => 
                           n11817, A => n9498, ZN => n9497);
   U9118 : OAI222_X1 port map( A1 => n11813, A2 => n8699, B1 => n11809, B2 => 
                           n8443, C1 => n11805, C2 => n8315, ZN => n9498);
   U9119 : AOI221_X1 port map( B1 => n10708, B2 => n11821, C1 => n11124, C2 => 
                           n11817, A => n9481, ZN => n9480);
   U9120 : OAI222_X1 port map( A1 => n11813, A2 => n8698, B1 => n11809, B2 => 
                           n8442, C1 => n11805, C2 => n8314, ZN => n9481);
   U9121 : AOI221_X1 port map( B1 => n10709, B2 => n11822, C1 => n11125, C2 => 
                           n11818, A => n9464, ZN => n9463);
   U9122 : OAI222_X1 port map( A1 => n11814, A2 => n8697, B1 => n11810, B2 => 
                           n8441, C1 => n11806, C2 => n8313, ZN => n9464);
   U9123 : AOI221_X1 port map( B1 => n10710, B2 => n11822, C1 => n11126, C2 => 
                           n11818, A => n9447, ZN => n9446);
   U9124 : OAI222_X1 port map( A1 => n11814, A2 => n8696, B1 => n11810, B2 => 
                           n8440, C1 => n11806, C2 => n8312, ZN => n9447);
   U9125 : AOI221_X1 port map( B1 => n10711, B2 => n11822, C1 => n11127, C2 => 
                           n11818, A => n9430, ZN => n9429);
   U9126 : OAI222_X1 port map( A1 => n11814, A2 => n8695, B1 => n11810, B2 => 
                           n8439, C1 => n11806, C2 => n8311, ZN => n9430);
   U9127 : AOI221_X1 port map( B1 => n10712, B2 => n11822, C1 => n11128, C2 => 
                           n11818, A => n9413, ZN => n9412);
   U9128 : OAI222_X1 port map( A1 => n11814, A2 => n8694, B1 => n11810, B2 => 
                           n8438, C1 => n11806, C2 => n8310, ZN => n9413);
   U9129 : AOI221_X1 port map( B1 => n10713, B2 => n11822, C1 => n11129, C2 => 
                           n11818, A => n9396, ZN => n9395);
   U9130 : OAI222_X1 port map( A1 => n11814, A2 => n8693, B1 => n11810, B2 => 
                           n8437, C1 => n11806, C2 => n8309, ZN => n9396);
   U9131 : AOI221_X1 port map( B1 => n10714, B2 => n11822, C1 => n11130, C2 => 
                           n11818, A => n9379, ZN => n9378);
   U9132 : OAI222_X1 port map( A1 => n11814, A2 => n8692, B1 => n11810, B2 => 
                           n8436, C1 => n11806, C2 => n8308, ZN => n9379);
   U9133 : AOI221_X1 port map( B1 => n10715, B2 => n11822, C1 => n11131, C2 => 
                           n11818, A => n9362, ZN => n9361);
   U9134 : OAI222_X1 port map( A1 => n11814, A2 => n8691, B1 => n11810, B2 => 
                           n8435, C1 => n11806, C2 => n8307, ZN => n9362);
   U9135 : AOI221_X1 port map( B1 => n10716, B2 => n11822, C1 => n11132, C2 => 
                           n11818, A => n9329, ZN => n9326);
   U9136 : OAI222_X1 port map( A1 => n11814, A2 => n8690, B1 => n11810, B2 => 
                           n8434, C1 => n11806, C2 => n8306, ZN => n9329);
   U9137 : AOI221_X1 port map( B1 => n11836, B2 => n9875, C1 => n11831, C2 => 
                           Out1_0_port, A => n9876, ZN => n9859);
   U9138 : OAI22_X1 port map( A1 => n11827, A2 => n8817, B1 => n11823, B2 => 
                           n9265, ZN => n9876);
   U9139 : NAND4_X1 port map( A1 => n9877, A2 => n9878, A3 => n9879, A4 => 
                           n9880, ZN => n9875);
   U9140 : AOI221_X1 port map( B1 => n10845, B2 => n11764, C1 => n10717, C2 => 
                           n11760, A => n9887, ZN => n9877);
   U9141 : AOI221_X1 port map( B1 => n11837, B2 => n9849, C1 => n11831, C2 => 
                           Out1_1_port, A => n9850, ZN => n9842);
   U9142 : OAI22_X1 port map( A1 => n11827, A2 => n8816, B1 => n11823, B2 => 
                           n9264, ZN => n9850);
   U9143 : NAND4_X1 port map( A1 => n9851, A2 => n9852, A3 => n9853, A4 => 
                           n9854, ZN => n9849);
   U9144 : AOI221_X1 port map( B1 => n10846, B2 => n11764, C1 => n10718, C2 => 
                           n11760, A => n9858, ZN => n9851);
   U9145 : AOI221_X1 port map( B1 => n11837, B2 => n9832, C1 => n11831, C2 => 
                           Out1_2_port, A => n9833, ZN => n9825);
   U9146 : OAI22_X1 port map( A1 => n11827, A2 => n8815, B1 => n11823, B2 => 
                           n9263, ZN => n9833);
   U9147 : NAND4_X1 port map( A1 => n9834, A2 => n9835, A3 => n9836, A4 => 
                           n9837, ZN => n9832);
   U9148 : AOI221_X1 port map( B1 => n10847, B2 => n11764, C1 => n10719, C2 => 
                           n11760, A => n9841, ZN => n9834);
   U9149 : AOI221_X1 port map( B1 => n11837, B2 => n9815, C1 => n11831, C2 => 
                           Out1_3_port, A => n9816, ZN => n9808);
   U9150 : OAI22_X1 port map( A1 => n11827, A2 => n8814, B1 => n11823, B2 => 
                           n9262, ZN => n9816);
   U9151 : NAND4_X1 port map( A1 => n9817, A2 => n9818, A3 => n9819, A4 => 
                           n9820, ZN => n9815);
   U9152 : AOI221_X1 port map( B1 => n10848, B2 => n11764, C1 => n10720, C2 => 
                           n11760, A => n9824, ZN => n9817);
   U9153 : AOI221_X1 port map( B1 => n11837, B2 => n9798, C1 => n11831, C2 => 
                           Out1_4_port, A => n9799, ZN => n9791);
   U9154 : OAI22_X1 port map( A1 => n11827, A2 => n8813, B1 => n11823, B2 => 
                           n9261, ZN => n9799);
   U9155 : NAND4_X1 port map( A1 => n9800, A2 => n9801, A3 => n9802, A4 => 
                           n9803, ZN => n9798);
   U9156 : AOI221_X1 port map( B1 => n10849, B2 => n11764, C1 => n10721, C2 => 
                           n11760, A => n9807, ZN => n9800);
   U9157 : AOI221_X1 port map( B1 => n11837, B2 => n9781, C1 => n11831, C2 => 
                           Out1_5_port, A => n9782, ZN => n9774);
   U9158 : OAI22_X1 port map( A1 => n11827, A2 => n8812, B1 => n11823, B2 => 
                           n9260, ZN => n9782);
   U9159 : NAND4_X1 port map( A1 => n9783, A2 => n9784, A3 => n9785, A4 => 
                           n9786, ZN => n9781);
   U9160 : AOI221_X1 port map( B1 => n10850, B2 => n11764, C1 => n10722, C2 => 
                           n11760, A => n9790, ZN => n9783);
   U9161 : AOI221_X1 port map( B1 => n11837, B2 => n9764, C1 => n11831, C2 => 
                           Out1_6_port, A => n9765, ZN => n9757);
   U9162 : OAI22_X1 port map( A1 => n11827, A2 => n8811, B1 => n11823, B2 => 
                           n9259, ZN => n9765);
   U9163 : NAND4_X1 port map( A1 => n9766, A2 => n9767, A3 => n9768, A4 => 
                           n9769, ZN => n9764);
   U9164 : AOI221_X1 port map( B1 => n10851, B2 => n11764, C1 => n10723, C2 => 
                           n11760, A => n9773, ZN => n9766);
   U9165 : AOI221_X1 port map( B1 => n11837, B2 => n9747, C1 => n11831, C2 => 
                           Out1_7_port, A => n9748, ZN => n9740);
   U9166 : OAI22_X1 port map( A1 => n11827, A2 => n8810, B1 => n11823, B2 => 
                           n9258, ZN => n9748);
   U9167 : NAND4_X1 port map( A1 => n9749, A2 => n9750, A3 => n9751, A4 => 
                           n9752, ZN => n9747);
   U9168 : AOI221_X1 port map( B1 => n10852, B2 => n11764, C1 => n10724, C2 => 
                           n11760, A => n9756, ZN => n9749);
   U9169 : AOI221_X1 port map( B1 => n11837, B2 => n9730, C1 => n11831, C2 => 
                           Out1_8_port, A => n9731, ZN => n9723);
   U9170 : OAI22_X1 port map( A1 => n11827, A2 => n8809, B1 => n11823, B2 => 
                           n9257, ZN => n9731);
   U9171 : NAND4_X1 port map( A1 => n9732, A2 => n9733, A3 => n9734, A4 => 
                           n9735, ZN => n9730);
   U9172 : AOI221_X1 port map( B1 => n10853, B2 => n11764, C1 => n10725, C2 => 
                           n11760, A => n9739, ZN => n9732);
   U9173 : AOI221_X1 port map( B1 => n11836, B2 => n9713, C1 => n11831, C2 => 
                           Out1_9_port, A => n9714, ZN => n9706);
   U9174 : OAI22_X1 port map( A1 => n11827, A2 => n8808, B1 => n11823, B2 => 
                           n9256, ZN => n9714);
   U9175 : NAND4_X1 port map( A1 => n9715, A2 => n9716, A3 => n9717, A4 => 
                           n9718, ZN => n9713);
   U9176 : AOI221_X1 port map( B1 => n10854, B2 => n11764, C1 => n10726, C2 => 
                           n11760, A => n9722, ZN => n9715);
   U9177 : AOI221_X1 port map( B1 => n11836, B2 => n9696, C1 => n11831, C2 => 
                           Out1_10_port, A => n9697, ZN => n9689);
   U9178 : OAI22_X1 port map( A1 => n11827, A2 => n8807, B1 => n11823, B2 => 
                           n9255, ZN => n9697);
   U9179 : NAND4_X1 port map( A1 => n9698, A2 => n9699, A3 => n9700, A4 => 
                           n9701, ZN => n9696);
   U9180 : AOI221_X1 port map( B1 => n10855, B2 => n11764, C1 => n10727, C2 => 
                           n11760, A => n9705, ZN => n9698);
   U9181 : AOI221_X1 port map( B1 => n11836, B2 => n9679, C1 => n11831, C2 => 
                           Out1_11_port, A => n9680, ZN => n9672);
   U9182 : OAI22_X1 port map( A1 => n11827, A2 => n8806, B1 => n11823, B2 => 
                           n9254, ZN => n9680);
   U9183 : NAND4_X1 port map( A1 => n9681, A2 => n9682, A3 => n9683, A4 => 
                           n9684, ZN => n9679);
   U9184 : AOI221_X1 port map( B1 => n10856, B2 => n11764, C1 => n10728, C2 => 
                           n11760, A => n9688, ZN => n9681);
   U9185 : AOI221_X1 port map( B1 => n11836, B2 => n9662, C1 => n11832, C2 => 
                           Out1_12_port, A => n9663, ZN => n9655);
   U9186 : OAI22_X1 port map( A1 => n11828, A2 => n8805, B1 => n11824, B2 => 
                           n9253, ZN => n9663);
   U9187 : NAND4_X1 port map( A1 => n9664, A2 => n9665, A3 => n9666, A4 => 
                           n9667, ZN => n9662);
   U9188 : AOI221_X1 port map( B1 => n10857, B2 => n11765, C1 => n10729, C2 => 
                           n11761, A => n9671, ZN => n9664);
   U9189 : AOI221_X1 port map( B1 => n11836, B2 => n9645, C1 => n11832, C2 => 
                           Out1_13_port, A => n9646, ZN => n9638);
   U9190 : OAI22_X1 port map( A1 => n11828, A2 => n8804, B1 => n11824, B2 => 
                           n9252, ZN => n9646);
   U9191 : NAND4_X1 port map( A1 => n9647, A2 => n9648, A3 => n9649, A4 => 
                           n9650, ZN => n9645);
   U9192 : AOI221_X1 port map( B1 => n10858, B2 => n11765, C1 => n10730, C2 => 
                           n11761, A => n9654, ZN => n9647);
   U9193 : AOI221_X1 port map( B1 => n11836, B2 => n9628, C1 => n11832, C2 => 
                           Out1_14_port, A => n9629, ZN => n9621);
   U9194 : OAI22_X1 port map( A1 => n11828, A2 => n8803, B1 => n11824, B2 => 
                           n9251, ZN => n9629);
   U9195 : NAND4_X1 port map( A1 => n9630, A2 => n9631, A3 => n9632, A4 => 
                           n9633, ZN => n9628);
   U9196 : AOI221_X1 port map( B1 => n10859, B2 => n11765, C1 => n10731, C2 => 
                           n11761, A => n9637, ZN => n9630);
   U9197 : AOI221_X1 port map( B1 => n11836, B2 => n9611, C1 => n11832, C2 => 
                           Out1_15_port, A => n9612, ZN => n9604);
   U9198 : OAI22_X1 port map( A1 => n11828, A2 => n8802, B1 => n11824, B2 => 
                           n9250, ZN => n9612);
   U9199 : NAND4_X1 port map( A1 => n9613, A2 => n9614, A3 => n9615, A4 => 
                           n9616, ZN => n9611);
   U9200 : AOI221_X1 port map( B1 => n10860, B2 => n11765, C1 => n10732, C2 => 
                           n11761, A => n9620, ZN => n9613);
   U9201 : AOI221_X1 port map( B1 => n11836, B2 => n9594, C1 => n11832, C2 => 
                           Out1_16_port, A => n9595, ZN => n9587);
   U9202 : OAI22_X1 port map( A1 => n11828, A2 => n8801, B1 => n11824, B2 => 
                           n9249, ZN => n9595);
   U9203 : NAND4_X1 port map( A1 => n9596, A2 => n9597, A3 => n9598, A4 => 
                           n9599, ZN => n9594);
   U9204 : AOI221_X1 port map( B1 => n10861, B2 => n11765, C1 => n10733, C2 => 
                           n11761, A => n9603, ZN => n9596);
   U9205 : AOI221_X1 port map( B1 => n11836, B2 => n9577, C1 => n11832, C2 => 
                           Out1_17_port, A => n9578, ZN => n9570);
   U9206 : OAI22_X1 port map( A1 => n11828, A2 => n8800, B1 => n11824, B2 => 
                           n9248, ZN => n9578);
   U9207 : NAND4_X1 port map( A1 => n9579, A2 => n9580, A3 => n9581, A4 => 
                           n9582, ZN => n9577);
   U9208 : AOI221_X1 port map( B1 => n10862, B2 => n11765, C1 => n10734, C2 => 
                           n11761, A => n9586, ZN => n9579);
   U9209 : AOI221_X1 port map( B1 => n11836, B2 => n9560, C1 => n11832, C2 => 
                           Out1_18_port, A => n9561, ZN => n9553);
   U9210 : OAI22_X1 port map( A1 => n11828, A2 => n8799, B1 => n11824, B2 => 
                           n9247, ZN => n9561);
   U9211 : NAND4_X1 port map( A1 => n9562, A2 => n9563, A3 => n9564, A4 => 
                           n9565, ZN => n9560);
   U9212 : AOI221_X1 port map( B1 => n10863, B2 => n11765, C1 => n10735, C2 => 
                           n11761, A => n9569, ZN => n9562);
   U9213 : AOI221_X1 port map( B1 => n11836, B2 => n9543, C1 => n11832, C2 => 
                           Out1_19_port, A => n9544, ZN => n9536);
   U9214 : OAI22_X1 port map( A1 => n11828, A2 => n8798, B1 => n11824, B2 => 
                           n9246, ZN => n9544);
   U9215 : NAND4_X1 port map( A1 => n9545, A2 => n9546, A3 => n9547, A4 => 
                           n9548, ZN => n9543);
   U9216 : AOI221_X1 port map( B1 => n10864, B2 => n11765, C1 => n10736, C2 => 
                           n11761, A => n9552, ZN => n9545);
   U9217 : AOI221_X1 port map( B1 => n11835, B2 => n9526, C1 => n11832, C2 => 
                           Out1_20_port, A => n9527, ZN => n9519);
   U9218 : OAI22_X1 port map( A1 => n11828, A2 => n8797, B1 => n11824, B2 => 
                           n9245, ZN => n9527);
   U9219 : NAND4_X1 port map( A1 => n9528, A2 => n9529, A3 => n9530, A4 => 
                           n9531, ZN => n9526);
   U9220 : AOI221_X1 port map( B1 => n10865, B2 => n11765, C1 => n10737, C2 => 
                           n11761, A => n9535, ZN => n9528);
   U9221 : AOI221_X1 port map( B1 => n11835, B2 => n9509, C1 => n11832, C2 => 
                           Out1_21_port, A => n9510, ZN => n9502);
   U9222 : OAI22_X1 port map( A1 => n11828, A2 => n8796, B1 => n11824, B2 => 
                           n9244, ZN => n9510);
   U9223 : NAND4_X1 port map( A1 => n9511, A2 => n9512, A3 => n9513, A4 => 
                           n9514, ZN => n9509);
   U9224 : AOI221_X1 port map( B1 => n10866, B2 => n11765, C1 => n10738, C2 => 
                           n11761, A => n9518, ZN => n9511);
   U9225 : AOI221_X1 port map( B1 => n11835, B2 => n9492, C1 => n11832, C2 => 
                           Out1_22_port, A => n9493, ZN => n9485);
   U9226 : OAI22_X1 port map( A1 => n11828, A2 => n8795, B1 => n11824, B2 => 
                           n9243, ZN => n9493);
   U9227 : NAND4_X1 port map( A1 => n9494, A2 => n9495, A3 => n9496, A4 => 
                           n9497, ZN => n9492);
   U9228 : AOI221_X1 port map( B1 => n10867, B2 => n11765, C1 => n10739, C2 => 
                           n11761, A => n9501, ZN => n9494);
   U9229 : AOI221_X1 port map( B1 => n11835, B2 => n9475, C1 => n11832, C2 => 
                           Out1_23_port, A => n9476, ZN => n9468);
   U9230 : OAI22_X1 port map( A1 => n11828, A2 => n8794, B1 => n11824, B2 => 
                           n9242, ZN => n9476);
   U9231 : NAND4_X1 port map( A1 => n9477, A2 => n9478, A3 => n9479, A4 => 
                           n9480, ZN => n9475);
   U9232 : AOI221_X1 port map( B1 => n10868, B2 => n11765, C1 => n10740, C2 => 
                           n11761, A => n9484, ZN => n9477);
   U9233 : AOI221_X1 port map( B1 => n11835, B2 => n9458, C1 => n11832, C2 => 
                           Out1_24_port, A => n9459, ZN => n9451);
   U9234 : OAI22_X1 port map( A1 => n11829, A2 => n8793, B1 => n11825, B2 => 
                           n9241, ZN => n9459);
   U9235 : NAND4_X1 port map( A1 => n9460, A2 => n9461, A3 => n9462, A4 => 
                           n9463, ZN => n9458);
   U9236 : AOI221_X1 port map( B1 => n10869, B2 => n11766, C1 => n10741, C2 => 
                           n11762, A => n9467, ZN => n9460);
   U9237 : AOI221_X1 port map( B1 => n11835, B2 => n9441, C1 => n11833, C2 => 
                           Out1_25_port, A => n9442, ZN => n9434);
   U9238 : OAI22_X1 port map( A1 => n11829, A2 => n8792, B1 => n11825, B2 => 
                           n9240, ZN => n9442);
   U9239 : NAND4_X1 port map( A1 => n9443, A2 => n9444, A3 => n9445, A4 => 
                           n9446, ZN => n9441);
   U9240 : AOI221_X1 port map( B1 => n10870, B2 => n11766, C1 => n10742, C2 => 
                           n11762, A => n9450, ZN => n9443);
   U9241 : AOI221_X1 port map( B1 => n11835, B2 => n9424, C1 => n11833, C2 => 
                           Out1_26_port, A => n9425, ZN => n9417);
   U9242 : OAI22_X1 port map( A1 => n11829, A2 => n8791, B1 => n11825, B2 => 
                           n9239, ZN => n9425);
   U9243 : NAND4_X1 port map( A1 => n9426, A2 => n9427, A3 => n9428, A4 => 
                           n9429, ZN => n9424);
   U9244 : AOI221_X1 port map( B1 => n10871, B2 => n11766, C1 => n10743, C2 => 
                           n11762, A => n9433, ZN => n9426);
   U9245 : AOI221_X1 port map( B1 => n11835, B2 => n9407, C1 => n11833, C2 => 
                           Out1_27_port, A => n9408, ZN => n9400);
   U9246 : OAI22_X1 port map( A1 => n11829, A2 => n8790, B1 => n11825, B2 => 
                           n9238, ZN => n9408);
   U9247 : NAND4_X1 port map( A1 => n9409, A2 => n9410, A3 => n9411, A4 => 
                           n9412, ZN => n9407);
   U9248 : AOI221_X1 port map( B1 => n10872, B2 => n11766, C1 => n10744, C2 => 
                           n11762, A => n9416, ZN => n9409);
   U9249 : AOI221_X1 port map( B1 => n11835, B2 => n9390, C1 => n11833, C2 => 
                           Out1_28_port, A => n9391, ZN => n9383);
   U9250 : OAI22_X1 port map( A1 => n11829, A2 => n8789, B1 => n11825, B2 => 
                           n9237, ZN => n9391);
   U9251 : NAND4_X1 port map( A1 => n9392, A2 => n9393, A3 => n9394, A4 => 
                           n9395, ZN => n9390);
   U9252 : AOI221_X1 port map( B1 => n10873, B2 => n11766, C1 => n10745, C2 => 
                           n11762, A => n9399, ZN => n9392);
   U9253 : AOI221_X1 port map( B1 => n11835, B2 => n9373, C1 => n11833, C2 => 
                           Out1_29_port, A => n9374, ZN => n9366);
   U9254 : OAI22_X1 port map( A1 => n11829, A2 => n8788, B1 => n11825, B2 => 
                           n9236, ZN => n9374);
   U9255 : NAND4_X1 port map( A1 => n9375, A2 => n9376, A3 => n9377, A4 => 
                           n9378, ZN => n9373);
   U9256 : AOI221_X1 port map( B1 => n10874, B2 => n11766, C1 => n10746, C2 => 
                           n11762, A => n9382, ZN => n9375);
   U9257 : AOI221_X1 port map( B1 => n11835, B2 => n9356, C1 => n11833, C2 => 
                           Out1_30_port, A => n9357, ZN => n9349);
   U9258 : OAI22_X1 port map( A1 => n11829, A2 => n8787, B1 => n11825, B2 => 
                           n9235, ZN => n9357);
   U9259 : NAND4_X1 port map( A1 => n9358, A2 => n9359, A3 => n9360, A4 => 
                           n9361, ZN => n9356);
   U9260 : AOI221_X1 port map( B1 => n10875, B2 => n11766, C1 => n10747, C2 => 
                           n11762, A => n9365, ZN => n9358);
   U9261 : AOI221_X1 port map( B1 => n11835, B2 => n9318, C1 => n11833, C2 => 
                           Out1_31_port, A => n9320, ZN => n9298);
   U9262 : OAI22_X1 port map( A1 => n11829, A2 => n8786, B1 => n11825, B2 => 
                           n9234, ZN => n9320);
   U9263 : NAND4_X1 port map( A1 => n9323, A2 => n9324, A3 => n9325, A4 => 
                           n9326, ZN => n9318);
   U9264 : AOI221_X1 port map( B1 => n10876, B2 => n11766, C1 => n10748, C2 => 
                           n11762, A => n9346, ZN => n9323);
   U9265 : NAND4_X1 port map( A1 => n9859, A2 => n9860, A3 => n9861, A4 => 
                           n9862, ZN => n7246);
   U9266 : AOI221_X1 port map( B1 => n7398, B2 => n11855, C1 => n7558, C2 => 
                           n11851, A => n9872, ZN => n9860);
   U9267 : AOI221_X1 port map( B1 => n7590, B2 => n11871, C1 => n10909, C2 => 
                           n11867, A => n9869, ZN => n9861);
   U9268 : AOI221_X1 port map( B1 => n7494, B2 => n11887, C1 => n10941, C2 => 
                           n11883, A => n9863, ZN => n9862);
   U9269 : NAND4_X1 port map( A1 => n9842, A2 => n9843, A3 => n9844, A4 => 
                           n9845, ZN => n7247);
   U9270 : AOI221_X1 port map( B1 => n7399, B2 => n11855, C1 => n7559, C2 => 
                           n11851, A => n9848, ZN => n9843);
   U9271 : AOI221_X1 port map( B1 => n7591, B2 => n11871, C1 => n10910, C2 => 
                           n11867, A => n9847, ZN => n9844);
   U9272 : AOI221_X1 port map( B1 => n7495, B2 => n11887, C1 => n10942, C2 => 
                           n11883, A => n9846, ZN => n9845);
   U9273 : NAND4_X1 port map( A1 => n9825, A2 => n9826, A3 => n9827, A4 => 
                           n9828, ZN => n7248);
   U9274 : AOI221_X1 port map( B1 => n7400, B2 => n11855, C1 => n7560, C2 => 
                           n11851, A => n9831, ZN => n9826);
   U9275 : AOI221_X1 port map( B1 => n7592, B2 => n11871, C1 => n10911, C2 => 
                           n11867, A => n9830, ZN => n9827);
   U9276 : AOI221_X1 port map( B1 => n7496, B2 => n11887, C1 => n10943, C2 => 
                           n11883, A => n9829, ZN => n9828);
   U9277 : NAND4_X1 port map( A1 => n9808, A2 => n9809, A3 => n9810, A4 => 
                           n9811, ZN => n7249);
   U9278 : AOI221_X1 port map( B1 => n7401, B2 => n11855, C1 => n7561, C2 => 
                           n11851, A => n9814, ZN => n9809);
   U9279 : AOI221_X1 port map( B1 => n7593, B2 => n11871, C1 => n10912, C2 => 
                           n11867, A => n9813, ZN => n9810);
   U9280 : AOI221_X1 port map( B1 => n7497, B2 => n11887, C1 => n10944, C2 => 
                           n11883, A => n9812, ZN => n9811);
   U9281 : NAND4_X1 port map( A1 => n9791, A2 => n9792, A3 => n9793, A4 => 
                           n9794, ZN => n7250);
   U9282 : AOI221_X1 port map( B1 => n7402, B2 => n11855, C1 => n7562, C2 => 
                           n11851, A => n9797, ZN => n9792);
   U9283 : AOI221_X1 port map( B1 => n7594, B2 => n11871, C1 => n10913, C2 => 
                           n11867, A => n9796, ZN => n9793);
   U9284 : AOI221_X1 port map( B1 => n7498, B2 => n11887, C1 => n10945, C2 => 
                           n11883, A => n9795, ZN => n9794);
   U9285 : NAND4_X1 port map( A1 => n9774, A2 => n9775, A3 => n9776, A4 => 
                           n9777, ZN => n7251);
   U9286 : AOI221_X1 port map( B1 => n7403, B2 => n11855, C1 => n7563, C2 => 
                           n11851, A => n9780, ZN => n9775);
   U9287 : AOI221_X1 port map( B1 => n7595, B2 => n11871, C1 => n10914, C2 => 
                           n11867, A => n9779, ZN => n9776);
   U9288 : AOI221_X1 port map( B1 => n7499, B2 => n11887, C1 => n10946, C2 => 
                           n11883, A => n9778, ZN => n9777);
   U9289 : NAND4_X1 port map( A1 => n9757, A2 => n9758, A3 => n9759, A4 => 
                           n9760, ZN => n7252);
   U9290 : AOI221_X1 port map( B1 => n7404, B2 => n11855, C1 => n7564, C2 => 
                           n11851, A => n9763, ZN => n9758);
   U9291 : AOI221_X1 port map( B1 => n7596, B2 => n11871, C1 => n10915, C2 => 
                           n11867, A => n9762, ZN => n9759);
   U9292 : AOI221_X1 port map( B1 => n7500, B2 => n11887, C1 => n10947, C2 => 
                           n11883, A => n9761, ZN => n9760);
   U9293 : NAND4_X1 port map( A1 => n9740, A2 => n9741, A3 => n9742, A4 => 
                           n9743, ZN => n7253);
   U9294 : AOI221_X1 port map( B1 => n7405, B2 => n11855, C1 => n7565, C2 => 
                           n11851, A => n9746, ZN => n9741);
   U9295 : AOI221_X1 port map( B1 => n7597, B2 => n11871, C1 => n10916, C2 => 
                           n11867, A => n9745, ZN => n9742);
   U9296 : AOI221_X1 port map( B1 => n7501, B2 => n11887, C1 => n10948, C2 => 
                           n11883, A => n9744, ZN => n9743);
   U9297 : NAND4_X1 port map( A1 => n9723, A2 => n9724, A3 => n9725, A4 => 
                           n9726, ZN => n7254);
   U9298 : AOI221_X1 port map( B1 => n7397, B2 => n11855, C1 => n7557, C2 => 
                           n11851, A => n9729, ZN => n9724);
   U9299 : AOI221_X1 port map( B1 => n7589, B2 => n11871, C1 => n10917, C2 => 
                           n11867, A => n9728, ZN => n9725);
   U9300 : AOI221_X1 port map( B1 => n7493, B2 => n11887, C1 => n10949, C2 => 
                           n11883, A => n9727, ZN => n9726);
   U9301 : NAND4_X1 port map( A1 => n9706, A2 => n9707, A3 => n9708, A4 => 
                           n9709, ZN => n7255);
   U9302 : AOI221_X1 port map( B1 => n7374, B2 => n11855, C1 => n7534, C2 => 
                           n11851, A => n9712, ZN => n9707);
   U9303 : AOI221_X1 port map( B1 => n7566, B2 => n11871, C1 => n10918, C2 => 
                           n11867, A => n9711, ZN => n9708);
   U9304 : AOI221_X1 port map( B1 => n7470, B2 => n11887, C1 => n10950, C2 => 
                           n11883, A => n9710, ZN => n9709);
   U9305 : NAND4_X1 port map( A1 => n9689, A2 => n9690, A3 => n9691, A4 => 
                           n9692, ZN => n7256);
   U9306 : AOI221_X1 port map( B1 => n7375, B2 => n11855, C1 => n7535, C2 => 
                           n11851, A => n9695, ZN => n9690);
   U9307 : AOI221_X1 port map( B1 => n7567, B2 => n11871, C1 => n10919, C2 => 
                           n11867, A => n9694, ZN => n9691);
   U9308 : AOI221_X1 port map( B1 => n7471, B2 => n11887, C1 => n10951, C2 => 
                           n11883, A => n9693, ZN => n9692);
   U9309 : NAND4_X1 port map( A1 => n9672, A2 => n9673, A3 => n9674, A4 => 
                           n9675, ZN => n7257);
   U9310 : AOI221_X1 port map( B1 => n7376, B2 => n11855, C1 => n7536, C2 => 
                           n11851, A => n9678, ZN => n9673);
   U9311 : AOI221_X1 port map( B1 => n7568, B2 => n11871, C1 => n10920, C2 => 
                           n11867, A => n9677, ZN => n9674);
   U9312 : AOI221_X1 port map( B1 => n7472, B2 => n11887, C1 => n10952, C2 => 
                           n11883, A => n9676, ZN => n9675);
   U9313 : NAND4_X1 port map( A1 => n9655, A2 => n9656, A3 => n9657, A4 => 
                           n9658, ZN => n7258);
   U9314 : AOI221_X1 port map( B1 => n7377, B2 => n11856, C1 => n7537, C2 => 
                           n11852, A => n9661, ZN => n9656);
   U9315 : AOI221_X1 port map( B1 => n7569, B2 => n11872, C1 => n10921, C2 => 
                           n11868, A => n9660, ZN => n9657);
   U9316 : AOI221_X1 port map( B1 => n7473, B2 => n11888, C1 => n10953, C2 => 
                           n11884, A => n9659, ZN => n9658);
   U9317 : NAND4_X1 port map( A1 => n9638, A2 => n9639, A3 => n9640, A4 => 
                           n9641, ZN => n7259);
   U9318 : AOI221_X1 port map( B1 => n7378, B2 => n11856, C1 => n7538, C2 => 
                           n11852, A => n9644, ZN => n9639);
   U9319 : AOI221_X1 port map( B1 => n7570, B2 => n11872, C1 => n10922, C2 => 
                           n11868, A => n9643, ZN => n9640);
   U9320 : AOI221_X1 port map( B1 => n7474, B2 => n11888, C1 => n10954, C2 => 
                           n11884, A => n9642, ZN => n9641);
   U9321 : NAND4_X1 port map( A1 => n9621, A2 => n9622, A3 => n9623, A4 => 
                           n9624, ZN => n7260);
   U9322 : AOI221_X1 port map( B1 => n7379, B2 => n11856, C1 => n7539, C2 => 
                           n11852, A => n9627, ZN => n9622);
   U9323 : AOI221_X1 port map( B1 => n7571, B2 => n11872, C1 => n10923, C2 => 
                           n11868, A => n9626, ZN => n9623);
   U9324 : AOI221_X1 port map( B1 => n7475, B2 => n11888, C1 => n10955, C2 => 
                           n11884, A => n9625, ZN => n9624);
   U9325 : NAND4_X1 port map( A1 => n9604, A2 => n9605, A3 => n9606, A4 => 
                           n9607, ZN => n7261);
   U9326 : AOI221_X1 port map( B1 => n7380, B2 => n11856, C1 => n7540, C2 => 
                           n11852, A => n9610, ZN => n9605);
   U9327 : AOI221_X1 port map( B1 => n7572, B2 => n11872, C1 => n10924, C2 => 
                           n11868, A => n9609, ZN => n9606);
   U9328 : AOI221_X1 port map( B1 => n7476, B2 => n11888, C1 => n10956, C2 => 
                           n11884, A => n9608, ZN => n9607);
   U9329 : NAND4_X1 port map( A1 => n9587, A2 => n9588, A3 => n9589, A4 => 
                           n9590, ZN => n7262);
   U9330 : AOI221_X1 port map( B1 => n7381, B2 => n11856, C1 => n7541, C2 => 
                           n11852, A => n9593, ZN => n9588);
   U9331 : AOI221_X1 port map( B1 => n7573, B2 => n11872, C1 => n10925, C2 => 
                           n11868, A => n9592, ZN => n9589);
   U9332 : AOI221_X1 port map( B1 => n7477, B2 => n11888, C1 => n10957, C2 => 
                           n11884, A => n9591, ZN => n9590);
   U9333 : NAND4_X1 port map( A1 => n9570, A2 => n9571, A3 => n9572, A4 => 
                           n9573, ZN => n7263);
   U9334 : AOI221_X1 port map( B1 => n7382, B2 => n11856, C1 => n7542, C2 => 
                           n11852, A => n9576, ZN => n9571);
   U9335 : AOI221_X1 port map( B1 => n7574, B2 => n11872, C1 => n10926, C2 => 
                           n11868, A => n9575, ZN => n9572);
   U9336 : AOI221_X1 port map( B1 => n7478, B2 => n11888, C1 => n10958, C2 => 
                           n11884, A => n9574, ZN => n9573);
   U9337 : NAND4_X1 port map( A1 => n9553, A2 => n9554, A3 => n9555, A4 => 
                           n9556, ZN => n7264);
   U9338 : AOI221_X1 port map( B1 => n7383, B2 => n11856, C1 => n7543, C2 => 
                           n11852, A => n9559, ZN => n9554);
   U9339 : AOI221_X1 port map( B1 => n7575, B2 => n11872, C1 => n10927, C2 => 
                           n11868, A => n9558, ZN => n9555);
   U9340 : AOI221_X1 port map( B1 => n7479, B2 => n11888, C1 => n10959, C2 => 
                           n11884, A => n9557, ZN => n9556);
   U9341 : NAND4_X1 port map( A1 => n9536, A2 => n9537, A3 => n9538, A4 => 
                           n9539, ZN => n7265);
   U9342 : AOI221_X1 port map( B1 => n7384, B2 => n11856, C1 => n7544, C2 => 
                           n11852, A => n9542, ZN => n9537);
   U9343 : AOI221_X1 port map( B1 => n7576, B2 => n11872, C1 => n10928, C2 => 
                           n11868, A => n9541, ZN => n9538);
   U9344 : AOI221_X1 port map( B1 => n7480, B2 => n11888, C1 => n10960, C2 => 
                           n11884, A => n9540, ZN => n9539);
   U9345 : NAND4_X1 port map( A1 => n9519, A2 => n9520, A3 => n9521, A4 => 
                           n9522, ZN => n7266);
   U9346 : AOI221_X1 port map( B1 => n7385, B2 => n11856, C1 => n7545, C2 => 
                           n11852, A => n9525, ZN => n9520);
   U9347 : AOI221_X1 port map( B1 => n7577, B2 => n11872, C1 => n10929, C2 => 
                           n11868, A => n9524, ZN => n9521);
   U9348 : AOI221_X1 port map( B1 => n7481, B2 => n11888, C1 => n10961, C2 => 
                           n11884, A => n9523, ZN => n9522);
   U9349 : NAND4_X1 port map( A1 => n9502, A2 => n9503, A3 => n9504, A4 => 
                           n9505, ZN => n7267);
   U9350 : AOI221_X1 port map( B1 => n7386, B2 => n11856, C1 => n7546, C2 => 
                           n11852, A => n9508, ZN => n9503);
   U9351 : AOI221_X1 port map( B1 => n7578, B2 => n11872, C1 => n10930, C2 => 
                           n11868, A => n9507, ZN => n9504);
   U9352 : AOI221_X1 port map( B1 => n7482, B2 => n11888, C1 => n10962, C2 => 
                           n11884, A => n9506, ZN => n9505);
   U9353 : NAND4_X1 port map( A1 => n9485, A2 => n9486, A3 => n9487, A4 => 
                           n9488, ZN => n7268);
   U9354 : AOI221_X1 port map( B1 => n7387, B2 => n11856, C1 => n7547, C2 => 
                           n11852, A => n9491, ZN => n9486);
   U9355 : AOI221_X1 port map( B1 => n7579, B2 => n11872, C1 => n10931, C2 => 
                           n11868, A => n9490, ZN => n9487);
   U9356 : AOI221_X1 port map( B1 => n7483, B2 => n11888, C1 => n10963, C2 => 
                           n11884, A => n9489, ZN => n9488);
   U9357 : NAND4_X1 port map( A1 => n9468, A2 => n9469, A3 => n9470, A4 => 
                           n9471, ZN => n7269);
   U9358 : AOI221_X1 port map( B1 => n7388, B2 => n11856, C1 => n7548, C2 => 
                           n11852, A => n9474, ZN => n9469);
   U9359 : AOI221_X1 port map( B1 => n7580, B2 => n11872, C1 => n10932, C2 => 
                           n11868, A => n9473, ZN => n9470);
   U9360 : AOI221_X1 port map( B1 => n7484, B2 => n11888, C1 => n10964, C2 => 
                           n11884, A => n9472, ZN => n9471);
   U9361 : NAND4_X1 port map( A1 => n9451, A2 => n9452, A3 => n9453, A4 => 
                           n9454, ZN => n7270);
   U9362 : AOI221_X1 port map( B1 => n7389, B2 => n11857, C1 => n7549, C2 => 
                           n11853, A => n9457, ZN => n9452);
   U9363 : AOI221_X1 port map( B1 => n7581, B2 => n11873, C1 => n10933, C2 => 
                           n11869, A => n9456, ZN => n9453);
   U9364 : AOI221_X1 port map( B1 => n7485, B2 => n11889, C1 => n10965, C2 => 
                           n11885, A => n9455, ZN => n9454);
   U9365 : NAND4_X1 port map( A1 => n9434, A2 => n9435, A3 => n9436, A4 => 
                           n9437, ZN => n7271);
   U9366 : AOI221_X1 port map( B1 => n7390, B2 => n11857, C1 => n7550, C2 => 
                           n11853, A => n9440, ZN => n9435);
   U9367 : AOI221_X1 port map( B1 => n7582, B2 => n11873, C1 => n10934, C2 => 
                           n11869, A => n9439, ZN => n9436);
   U9368 : AOI221_X1 port map( B1 => n7486, B2 => n11889, C1 => n10966, C2 => 
                           n11885, A => n9438, ZN => n9437);
   U9369 : NAND4_X1 port map( A1 => n9417, A2 => n9418, A3 => n9419, A4 => 
                           n9420, ZN => n7272);
   U9370 : AOI221_X1 port map( B1 => n7391, B2 => n11857, C1 => n7551, C2 => 
                           n11853, A => n9423, ZN => n9418);
   U9371 : AOI221_X1 port map( B1 => n7583, B2 => n11873, C1 => n10935, C2 => 
                           n11869, A => n9422, ZN => n9419);
   U9372 : AOI221_X1 port map( B1 => n7487, B2 => n11889, C1 => n10967, C2 => 
                           n11885, A => n9421, ZN => n9420);
   U9373 : NAND4_X1 port map( A1 => n9400, A2 => n9401, A3 => n9402, A4 => 
                           n9403, ZN => n7273);
   U9374 : AOI221_X1 port map( B1 => n7392, B2 => n11857, C1 => n7552, C2 => 
                           n11853, A => n9406, ZN => n9401);
   U9375 : AOI221_X1 port map( B1 => n7584, B2 => n11873, C1 => n10936, C2 => 
                           n11869, A => n9405, ZN => n9402);
   U9376 : AOI221_X1 port map( B1 => n7488, B2 => n11889, C1 => n10968, C2 => 
                           n11885, A => n9404, ZN => n9403);
   U9377 : NAND4_X1 port map( A1 => n9383, A2 => n9384, A3 => n9385, A4 => 
                           n9386, ZN => n7274);
   U9378 : AOI221_X1 port map( B1 => n7393, B2 => n11857, C1 => n7553, C2 => 
                           n11853, A => n9389, ZN => n9384);
   U9379 : AOI221_X1 port map( B1 => n7585, B2 => n11873, C1 => n10937, C2 => 
                           n11869, A => n9388, ZN => n9385);
   U9380 : AOI221_X1 port map( B1 => n7489, B2 => n11889, C1 => n10969, C2 => 
                           n11885, A => n9387, ZN => n9386);
   U9381 : NAND4_X1 port map( A1 => n9366, A2 => n9367, A3 => n9368, A4 => 
                           n9369, ZN => n7275);
   U9382 : AOI221_X1 port map( B1 => n7394, B2 => n11857, C1 => n7554, C2 => 
                           n11853, A => n9372, ZN => n9367);
   U9383 : AOI221_X1 port map( B1 => n7586, B2 => n11873, C1 => n10938, C2 => 
                           n11869, A => n9371, ZN => n9368);
   U9384 : AOI221_X1 port map( B1 => n7490, B2 => n11889, C1 => n10970, C2 => 
                           n11885, A => n9370, ZN => n9369);
   U9385 : NAND4_X1 port map( A1 => n9349, A2 => n9350, A3 => n9351, A4 => 
                           n9352, ZN => n7276);
   U9386 : AOI221_X1 port map( B1 => n7395, B2 => n11857, C1 => n7555, C2 => 
                           n11853, A => n9355, ZN => n9350);
   U9387 : AOI221_X1 port map( B1 => n7587, B2 => n11873, C1 => n10939, C2 => 
                           n11869, A => n9354, ZN => n9351);
   U9388 : AOI221_X1 port map( B1 => n7491, B2 => n11889, C1 => n10971, C2 => 
                           n11885, A => n9353, ZN => n9352);
   U9389 : NAND4_X1 port map( A1 => n9298, A2 => n9299, A3 => n9300, A4 => 
                           n9301, ZN => n7277);
   U9390 : AOI221_X1 port map( B1 => n7396, B2 => n11857, C1 => n7556, C2 => 
                           n11853, A => n9314, ZN => n9299);
   U9391 : AOI221_X1 port map( B1 => n7588, B2 => n11873, C1 => n10940, C2 => 
                           n11869, A => n9309, ZN => n9300);
   U9392 : AOI221_X1 port map( B1 => n7492, B2 => n11889, C1 => n10972, C2 => 
                           n11885, A => n9304, ZN => n9301);
   U9393 : AOI221_X1 port map( B1 => n11681, B2 => n10685, C1 => n11677, C2 => 
                           n11101, A => n10471, ZN => n10470);
   U9394 : OAI222_X1 port map( A1 => n8721, A2 => n11673, B1 => n8465, B2 => 
                           n11669, C1 => n8337, C2 => n11665, ZN => n10471);
   U9395 : AOI221_X1 port map( B1 => n11681, B2 => n10686, C1 => n11677, C2 => 
                           n11102, A => n10445, ZN => n10444);
   U9396 : OAI222_X1 port map( A1 => n8720, A2 => n11673, B1 => n8464, B2 => 
                           n11669, C1 => n8336, C2 => n11665, ZN => n10445);
   U9397 : AOI221_X1 port map( B1 => n11681, B2 => n10687, C1 => n11677, C2 => 
                           n11103, A => n10428, ZN => n10427);
   U9398 : OAI222_X1 port map( A1 => n8719, A2 => n11673, B1 => n8463, B2 => 
                           n11669, C1 => n8335, C2 => n11665, ZN => n10428);
   U9399 : AOI221_X1 port map( B1 => n11681, B2 => n10688, C1 => n11677, C2 => 
                           n11104, A => n10411, ZN => n10410);
   U9400 : OAI222_X1 port map( A1 => n8718, A2 => n11673, B1 => n8462, B2 => 
                           n11669, C1 => n8334, C2 => n11665, ZN => n10411);
   U9401 : AOI221_X1 port map( B1 => n11681, B2 => n10689, C1 => n11677, C2 => 
                           n11105, A => n10394, ZN => n10393);
   U9402 : OAI222_X1 port map( A1 => n8717, A2 => n11673, B1 => n8461, B2 => 
                           n11669, C1 => n8333, C2 => n11665, ZN => n10394);
   U9403 : AOI221_X1 port map( B1 => n11681, B2 => n10690, C1 => n11677, C2 => 
                           n11106, A => n10377, ZN => n10376);
   U9404 : OAI222_X1 port map( A1 => n8716, A2 => n11673, B1 => n8460, B2 => 
                           n11669, C1 => n8332, C2 => n11665, ZN => n10377);
   U9405 : AOI221_X1 port map( B1 => n11681, B2 => n10691, C1 => n11677, C2 => 
                           n11107, A => n10360, ZN => n10359);
   U9406 : OAI222_X1 port map( A1 => n8715, A2 => n11673, B1 => n8459, B2 => 
                           n11669, C1 => n8331, C2 => n11665, ZN => n10360);
   U9407 : AOI221_X1 port map( B1 => n11681, B2 => n10692, C1 => n11677, C2 => 
                           n11108, A => n10343, ZN => n10342);
   U9408 : OAI222_X1 port map( A1 => n8714, A2 => n11673, B1 => n8458, B2 => 
                           n11669, C1 => n8330, C2 => n11665, ZN => n10343);
   U9409 : AOI221_X1 port map( B1 => n11681, B2 => n10693, C1 => n11677, C2 => 
                           n11109, A => n10326, ZN => n10325);
   U9410 : OAI222_X1 port map( A1 => n8713, A2 => n11673, B1 => n8457, B2 => 
                           n11669, C1 => n8329, C2 => n11665, ZN => n10326);
   U9411 : AOI221_X1 port map( B1 => n11681, B2 => n10694, C1 => n11677, C2 => 
                           n11110, A => n10309, ZN => n10308);
   U9412 : OAI222_X1 port map( A1 => n8712, A2 => n11673, B1 => n8456, B2 => 
                           n11669, C1 => n8328, C2 => n11665, ZN => n10309);
   U9413 : AOI221_X1 port map( B1 => n11681, B2 => n10695, C1 => n11677, C2 => 
                           n11111, A => n10292, ZN => n10291);
   U9414 : OAI222_X1 port map( A1 => n8711, A2 => n11673, B1 => n8455, B2 => 
                           n11669, C1 => n8327, C2 => n11665, ZN => n10292);
   U9415 : AOI221_X1 port map( B1 => n11681, B2 => n10696, C1 => n11677, C2 => 
                           n11112, A => n10275, ZN => n10274);
   U9416 : OAI222_X1 port map( A1 => n8710, A2 => n11673, B1 => n8454, B2 => 
                           n11669, C1 => n8326, C2 => n11665, ZN => n10275);
   U9417 : AOI221_X1 port map( B1 => n11682, B2 => n10697, C1 => n11678, C2 => 
                           n11113, A => n10258, ZN => n10257);
   U9418 : OAI222_X1 port map( A1 => n8709, A2 => n11674, B1 => n8453, B2 => 
                           n11670, C1 => n8325, C2 => n11666, ZN => n10258);
   U9419 : AOI221_X1 port map( B1 => n11682, B2 => n10698, C1 => n11678, C2 => 
                           n11114, A => n10241, ZN => n10240);
   U9420 : OAI222_X1 port map( A1 => n8708, A2 => n11674, B1 => n8452, B2 => 
                           n11670, C1 => n8324, C2 => n11666, ZN => n10241);
   U9421 : AOI221_X1 port map( B1 => n11682, B2 => n10699, C1 => n11678, C2 => 
                           n11115, A => n10224, ZN => n10223);
   U9422 : OAI222_X1 port map( A1 => n8707, A2 => n11674, B1 => n8451, B2 => 
                           n11670, C1 => n8323, C2 => n11666, ZN => n10224);
   U9423 : AOI221_X1 port map( B1 => n11682, B2 => n10700, C1 => n11678, C2 => 
                           n11116, A => n10207, ZN => n10206);
   U9424 : OAI222_X1 port map( A1 => n8706, A2 => n11674, B1 => n8450, B2 => 
                           n11670, C1 => n8322, C2 => n11666, ZN => n10207);
   U9425 : AOI221_X1 port map( B1 => n11682, B2 => n10701, C1 => n11678, C2 => 
                           n11117, A => n10190, ZN => n10189);
   U9426 : OAI222_X1 port map( A1 => n8705, A2 => n11674, B1 => n8449, B2 => 
                           n11670, C1 => n8321, C2 => n11666, ZN => n10190);
   U9427 : AOI221_X1 port map( B1 => n11682, B2 => n10702, C1 => n11678, C2 => 
                           n11118, A => n10173, ZN => n10172);
   U9428 : OAI222_X1 port map( A1 => n8704, A2 => n11674, B1 => n8448, B2 => 
                           n11670, C1 => n8320, C2 => n11666, ZN => n10173);
   U9429 : AOI221_X1 port map( B1 => n11682, B2 => n10703, C1 => n11678, C2 => 
                           n11119, A => n10156, ZN => n10155);
   U9430 : OAI222_X1 port map( A1 => n8703, A2 => n11674, B1 => n8447, B2 => 
                           n11670, C1 => n8319, C2 => n11666, ZN => n10156);
   U9431 : AOI221_X1 port map( B1 => n11682, B2 => n10704, C1 => n11678, C2 => 
                           n11120, A => n10139, ZN => n10138);
   U9432 : OAI222_X1 port map( A1 => n8702, A2 => n11674, B1 => n8446, B2 => 
                           n11670, C1 => n8318, C2 => n11666, ZN => n10139);
   U9433 : AOI221_X1 port map( B1 => n11682, B2 => n10705, C1 => n11678, C2 => 
                           n11121, A => n10122, ZN => n10121);
   U9434 : OAI222_X1 port map( A1 => n8701, A2 => n11674, B1 => n8445, B2 => 
                           n11670, C1 => n8317, C2 => n11666, ZN => n10122);
   U9435 : AOI221_X1 port map( B1 => n11682, B2 => n10706, C1 => n11678, C2 => 
                           n11122, A => n10105, ZN => n10104);
   U9436 : OAI222_X1 port map( A1 => n8700, A2 => n11674, B1 => n8444, B2 => 
                           n11670, C1 => n8316, C2 => n11666, ZN => n10105);
   U9437 : AOI221_X1 port map( B1 => n11682, B2 => n10707, C1 => n11678, C2 => 
                           n11123, A => n10088, ZN => n10087);
   U9438 : OAI222_X1 port map( A1 => n8699, A2 => n11674, B1 => n8443, B2 => 
                           n11670, C1 => n8315, C2 => n11666, ZN => n10088);
   U9439 : AOI221_X1 port map( B1 => n11682, B2 => n10708, C1 => n11678, C2 => 
                           n11124, A => n10071, ZN => n10070);
   U9440 : OAI222_X1 port map( A1 => n8698, A2 => n11674, B1 => n8442, B2 => 
                           n11670, C1 => n8314, C2 => n11666, ZN => n10071);
   U9441 : AOI221_X1 port map( B1 => n11683, B2 => n10709, C1 => n11679, C2 => 
                           n11125, A => n10054, ZN => n10053);
   U9442 : OAI222_X1 port map( A1 => n8697, A2 => n11675, B1 => n8441, B2 => 
                           n11671, C1 => n8313, C2 => n11667, ZN => n10054);
   U9443 : AOI221_X1 port map( B1 => n11683, B2 => n10710, C1 => n11679, C2 => 
                           n11126, A => n10037, ZN => n10036);
   U9444 : OAI222_X1 port map( A1 => n8696, A2 => n11675, B1 => n8440, B2 => 
                           n11671, C1 => n8312, C2 => n11667, ZN => n10037);
   U9445 : AOI221_X1 port map( B1 => n11683, B2 => n10711, C1 => n11679, C2 => 
                           n11127, A => n10020, ZN => n10019);
   U9446 : OAI222_X1 port map( A1 => n8695, A2 => n11675, B1 => n8439, B2 => 
                           n11671, C1 => n8311, C2 => n11667, ZN => n10020);
   U9447 : AOI221_X1 port map( B1 => n11683, B2 => n10712, C1 => n11679, C2 => 
                           n11128, A => n10003, ZN => n10002);
   U9448 : OAI222_X1 port map( A1 => n8694, A2 => n11675, B1 => n8438, B2 => 
                           n11671, C1 => n8310, C2 => n11667, ZN => n10003);
   U9449 : AOI221_X1 port map( B1 => n11683, B2 => n10713, C1 => n11679, C2 => 
                           n11129, A => n9986, ZN => n9985);
   U9450 : OAI222_X1 port map( A1 => n8693, A2 => n11675, B1 => n8437, B2 => 
                           n11671, C1 => n8309, C2 => n11667, ZN => n9986);
   U9451 : AOI221_X1 port map( B1 => n11683, B2 => n10714, C1 => n11679, C2 => 
                           n11130, A => n9969, ZN => n9968);
   U9452 : OAI222_X1 port map( A1 => n8692, A2 => n11675, B1 => n8436, B2 => 
                           n11671, C1 => n8308, C2 => n11667, ZN => n9969);
   U9453 : AOI221_X1 port map( B1 => n11683, B2 => n10715, C1 => n11679, C2 => 
                           n11131, A => n9952, ZN => n9951);
   U9454 : OAI222_X1 port map( A1 => n8691, A2 => n11675, B1 => n8435, B2 => 
                           n11671, C1 => n8307, C2 => n11667, ZN => n9952);
   U9455 : AOI221_X1 port map( B1 => n11683, B2 => n10716, C1 => n11679, C2 => 
                           n11132, A => n9919, ZN => n9916);
   U9456 : OAI222_X1 port map( A1 => n8690, A2 => n11675, B1 => n8434, B2 => 
                           n11671, C1 => n8306, C2 => n11667, ZN => n9919);
   U9457 : AOI221_X1 port map( B1 => n11697, B2 => n10465, C1 => n11692, C2 => 
                           Out2_0_port, A => n10466, ZN => n10449);
   U9458 : OAI22_X1 port map( A1 => n8817, A2 => n11688, B1 => n9265, B2 => 
                           n11684, ZN => n10466);
   U9459 : NAND4_X1 port map( A1 => n10467, A2 => n10468, A3 => n10469, A4 => 
                           n10470, ZN => n10465);
   U9460 : AOI221_X1 port map( B1 => n11625, B2 => n10845, C1 => n11621, C2 => 
                           n10717, A => n10477, ZN => n10467);
   U9461 : AOI221_X1 port map( B1 => n11698, B2 => n10439, C1 => n11692, C2 => 
                           Out2_1_port, A => n10440, ZN => n10432);
   U9462 : OAI22_X1 port map( A1 => n8816, A2 => n11688, B1 => n9264, B2 => 
                           n11684, ZN => n10440);
   U9463 : NAND4_X1 port map( A1 => n10441, A2 => n10442, A3 => n10443, A4 => 
                           n10444, ZN => n10439);
   U9464 : AOI221_X1 port map( B1 => n11625, B2 => n10846, C1 => n11621, C2 => 
                           n10718, A => n10448, ZN => n10441);
   U9465 : AOI221_X1 port map( B1 => n11698, B2 => n10422, C1 => n11692, C2 => 
                           Out2_2_port, A => n10423, ZN => n10415);
   U9466 : OAI22_X1 port map( A1 => n8815, A2 => n11688, B1 => n9263, B2 => 
                           n11684, ZN => n10423);
   U9467 : NAND4_X1 port map( A1 => n10424, A2 => n10425, A3 => n10426, A4 => 
                           n10427, ZN => n10422);
   U9468 : AOI221_X1 port map( B1 => n11625, B2 => n10847, C1 => n11621, C2 => 
                           n10719, A => n10431, ZN => n10424);
   U9469 : AOI221_X1 port map( B1 => n11698, B2 => n10405, C1 => n11692, C2 => 
                           Out2_3_port, A => n10406, ZN => n10398);
   U9470 : OAI22_X1 port map( A1 => n8814, A2 => n11688, B1 => n9262, B2 => 
                           n11684, ZN => n10406);
   U9471 : NAND4_X1 port map( A1 => n10407, A2 => n10408, A3 => n10409, A4 => 
                           n10410, ZN => n10405);
   U9472 : AOI221_X1 port map( B1 => n11625, B2 => n10848, C1 => n11621, C2 => 
                           n10720, A => n10414, ZN => n10407);
   U9473 : AOI221_X1 port map( B1 => n11698, B2 => n10388, C1 => n11692, C2 => 
                           Out2_4_port, A => n10389, ZN => n10381);
   U9474 : OAI22_X1 port map( A1 => n8813, A2 => n11688, B1 => n9261, B2 => 
                           n11684, ZN => n10389);
   U9475 : NAND4_X1 port map( A1 => n10390, A2 => n10391, A3 => n10392, A4 => 
                           n10393, ZN => n10388);
   U9476 : AOI221_X1 port map( B1 => n11625, B2 => n10849, C1 => n11621, C2 => 
                           n10721, A => n10397, ZN => n10390);
   U9477 : AOI221_X1 port map( B1 => n11698, B2 => n10371, C1 => n11692, C2 => 
                           Out2_5_port, A => n10372, ZN => n10364);
   U9478 : OAI22_X1 port map( A1 => n8812, A2 => n11688, B1 => n9260, B2 => 
                           n11684, ZN => n10372);
   U9479 : NAND4_X1 port map( A1 => n10373, A2 => n10374, A3 => n10375, A4 => 
                           n10376, ZN => n10371);
   U9480 : AOI221_X1 port map( B1 => n11625, B2 => n10850, C1 => n11621, C2 => 
                           n10722, A => n10380, ZN => n10373);
   U9481 : AOI221_X1 port map( B1 => n11698, B2 => n10354, C1 => n11692, C2 => 
                           Out2_6_port, A => n10355, ZN => n10347);
   U9482 : OAI22_X1 port map( A1 => n8811, A2 => n11688, B1 => n9259, B2 => 
                           n11684, ZN => n10355);
   U9483 : NAND4_X1 port map( A1 => n10356, A2 => n10357, A3 => n10358, A4 => 
                           n10359, ZN => n10354);
   U9484 : AOI221_X1 port map( B1 => n11625, B2 => n10851, C1 => n11621, C2 => 
                           n10723, A => n10363, ZN => n10356);
   U9485 : AOI221_X1 port map( B1 => n11698, B2 => n10337, C1 => n11692, C2 => 
                           Out2_7_port, A => n10338, ZN => n10330);
   U9486 : OAI22_X1 port map( A1 => n8810, A2 => n11688, B1 => n9258, B2 => 
                           n11684, ZN => n10338);
   U9487 : NAND4_X1 port map( A1 => n10339, A2 => n10340, A3 => n10341, A4 => 
                           n10342, ZN => n10337);
   U9488 : AOI221_X1 port map( B1 => n11625, B2 => n10852, C1 => n11621, C2 => 
                           n10724, A => n10346, ZN => n10339);
   U9489 : AOI221_X1 port map( B1 => n11698, B2 => n10320, C1 => n11692, C2 => 
                           Out2_8_port, A => n10321, ZN => n10313);
   U9490 : OAI22_X1 port map( A1 => n8809, A2 => n11688, B1 => n9257, B2 => 
                           n11684, ZN => n10321);
   U9491 : NAND4_X1 port map( A1 => n10322, A2 => n10323, A3 => n10324, A4 => 
                           n10325, ZN => n10320);
   U9492 : AOI221_X1 port map( B1 => n11625, B2 => n10853, C1 => n11621, C2 => 
                           n10725, A => n10329, ZN => n10322);
   U9493 : AOI221_X1 port map( B1 => n11697, B2 => n10303, C1 => n11692, C2 => 
                           Out2_9_port, A => n10304, ZN => n10296);
   U9494 : OAI22_X1 port map( A1 => n8808, A2 => n11688, B1 => n9256, B2 => 
                           n11684, ZN => n10304);
   U9495 : NAND4_X1 port map( A1 => n10305, A2 => n10306, A3 => n10307, A4 => 
                           n10308, ZN => n10303);
   U9496 : AOI221_X1 port map( B1 => n11625, B2 => n10854, C1 => n11621, C2 => 
                           n10726, A => n10312, ZN => n10305);
   U9497 : AOI221_X1 port map( B1 => n11697, B2 => n10286, C1 => n11692, C2 => 
                           Out2_10_port, A => n10287, ZN => n10279);
   U9498 : OAI22_X1 port map( A1 => n8807, A2 => n11688, B1 => n9255, B2 => 
                           n11684, ZN => n10287);
   U9499 : NAND4_X1 port map( A1 => n10288, A2 => n10289, A3 => n10290, A4 => 
                           n10291, ZN => n10286);
   U9500 : AOI221_X1 port map( B1 => n11625, B2 => n10855, C1 => n11621, C2 => 
                           n10727, A => n10295, ZN => n10288);
   U9501 : AOI221_X1 port map( B1 => n11697, B2 => n10269, C1 => n11692, C2 => 
                           Out2_11_port, A => n10270, ZN => n10262);
   U9502 : OAI22_X1 port map( A1 => n8806, A2 => n11688, B1 => n9254, B2 => 
                           n11684, ZN => n10270);
   U9503 : NAND4_X1 port map( A1 => n10271, A2 => n10272, A3 => n10273, A4 => 
                           n10274, ZN => n10269);
   U9504 : AOI221_X1 port map( B1 => n11625, B2 => n10856, C1 => n11621, C2 => 
                           n10728, A => n10278, ZN => n10271);
   U9505 : AOI221_X1 port map( B1 => n11697, B2 => n10252, C1 => n11693, C2 => 
                           Out2_12_port, A => n10253, ZN => n10245);
   U9506 : OAI22_X1 port map( A1 => n8805, A2 => n11689, B1 => n9253, B2 => 
                           n11685, ZN => n10253);
   U9507 : NAND4_X1 port map( A1 => n10254, A2 => n10255, A3 => n10256, A4 => 
                           n10257, ZN => n10252);
   U9508 : AOI221_X1 port map( B1 => n11626, B2 => n10857, C1 => n11622, C2 => 
                           n10729, A => n10261, ZN => n10254);
   U9509 : AOI221_X1 port map( B1 => n11697, B2 => n10235, C1 => n11693, C2 => 
                           Out2_13_port, A => n10236, ZN => n10228);
   U9510 : OAI22_X1 port map( A1 => n8804, A2 => n11689, B1 => n9252, B2 => 
                           n11685, ZN => n10236);
   U9511 : NAND4_X1 port map( A1 => n10237, A2 => n10238, A3 => n10239, A4 => 
                           n10240, ZN => n10235);
   U9512 : AOI221_X1 port map( B1 => n11626, B2 => n10858, C1 => n11622, C2 => 
                           n10730, A => n10244, ZN => n10237);
   U9513 : AOI221_X1 port map( B1 => n11697, B2 => n10218, C1 => n11693, C2 => 
                           Out2_14_port, A => n10219, ZN => n10211);
   U9514 : OAI22_X1 port map( A1 => n8803, A2 => n11689, B1 => n9251, B2 => 
                           n11685, ZN => n10219);
   U9515 : NAND4_X1 port map( A1 => n10220, A2 => n10221, A3 => n10222, A4 => 
                           n10223, ZN => n10218);
   U9516 : AOI221_X1 port map( B1 => n11626, B2 => n10859, C1 => n11622, C2 => 
                           n10731, A => n10227, ZN => n10220);
   U9517 : AOI221_X1 port map( B1 => n11697, B2 => n10201, C1 => n11693, C2 => 
                           Out2_15_port, A => n10202, ZN => n10194);
   U9518 : OAI22_X1 port map( A1 => n8802, A2 => n11689, B1 => n9250, B2 => 
                           n11685, ZN => n10202);
   U9519 : NAND4_X1 port map( A1 => n10203, A2 => n10204, A3 => n10205, A4 => 
                           n10206, ZN => n10201);
   U9520 : AOI221_X1 port map( B1 => n11626, B2 => n10860, C1 => n11622, C2 => 
                           n10732, A => n10210, ZN => n10203);
   U9521 : AOI221_X1 port map( B1 => n11697, B2 => n10184, C1 => n11693, C2 => 
                           Out2_16_port, A => n10185, ZN => n10177);
   U9522 : OAI22_X1 port map( A1 => n8801, A2 => n11689, B1 => n9249, B2 => 
                           n11685, ZN => n10185);
   U9523 : NAND4_X1 port map( A1 => n10186, A2 => n10187, A3 => n10188, A4 => 
                           n10189, ZN => n10184);
   U9524 : AOI221_X1 port map( B1 => n11626, B2 => n10861, C1 => n11622, C2 => 
                           n10733, A => n10193, ZN => n10186);
   U9525 : AOI221_X1 port map( B1 => n11697, B2 => n10167, C1 => n11693, C2 => 
                           Out2_17_port, A => n10168, ZN => n10160);
   U9526 : OAI22_X1 port map( A1 => n8800, A2 => n11689, B1 => n9248, B2 => 
                           n11685, ZN => n10168);
   U9527 : NAND4_X1 port map( A1 => n10169, A2 => n10170, A3 => n10171, A4 => 
                           n10172, ZN => n10167);
   U9528 : AOI221_X1 port map( B1 => n11626, B2 => n10862, C1 => n11622, C2 => 
                           n10734, A => n10176, ZN => n10169);
   U9529 : AOI221_X1 port map( B1 => n11697, B2 => n10150, C1 => n11693, C2 => 
                           Out2_18_port, A => n10151, ZN => n10143);
   U9530 : OAI22_X1 port map( A1 => n8799, A2 => n11689, B1 => n9247, B2 => 
                           n11685, ZN => n10151);
   U9531 : NAND4_X1 port map( A1 => n10152, A2 => n10153, A3 => n10154, A4 => 
                           n10155, ZN => n10150);
   U9532 : AOI221_X1 port map( B1 => n11626, B2 => n10863, C1 => n11622, C2 => 
                           n10735, A => n10159, ZN => n10152);
   U9533 : AOI221_X1 port map( B1 => n11697, B2 => n10133, C1 => n11693, C2 => 
                           Out2_19_port, A => n10134, ZN => n10126);
   U9534 : OAI22_X1 port map( A1 => n8798, A2 => n11689, B1 => n9246, B2 => 
                           n11685, ZN => n10134);
   U9535 : NAND4_X1 port map( A1 => n10135, A2 => n10136, A3 => n10137, A4 => 
                           n10138, ZN => n10133);
   U9536 : AOI221_X1 port map( B1 => n11626, B2 => n10864, C1 => n11622, C2 => 
                           n10736, A => n10142, ZN => n10135);
   U9537 : AOI221_X1 port map( B1 => n11696, B2 => n10116, C1 => n11693, C2 => 
                           Out2_20_port, A => n10117, ZN => n10109);
   U9538 : OAI22_X1 port map( A1 => n8797, A2 => n11689, B1 => n9245, B2 => 
                           n11685, ZN => n10117);
   U9539 : NAND4_X1 port map( A1 => n10118, A2 => n10119, A3 => n10120, A4 => 
                           n10121, ZN => n10116);
   U9540 : AOI221_X1 port map( B1 => n11626, B2 => n10865, C1 => n11622, C2 => 
                           n10737, A => n10125, ZN => n10118);
   U9541 : AOI221_X1 port map( B1 => n11696, B2 => n10099, C1 => n11693, C2 => 
                           Out2_21_port, A => n10100, ZN => n10092);
   U9542 : OAI22_X1 port map( A1 => n8796, A2 => n11689, B1 => n9244, B2 => 
                           n11685, ZN => n10100);
   U9543 : NAND4_X1 port map( A1 => n10101, A2 => n10102, A3 => n10103, A4 => 
                           n10104, ZN => n10099);
   U9544 : AOI221_X1 port map( B1 => n11626, B2 => n10866, C1 => n11622, C2 => 
                           n10738, A => n10108, ZN => n10101);
   U9545 : AOI221_X1 port map( B1 => n11696, B2 => n10082, C1 => n11693, C2 => 
                           Out2_22_port, A => n10083, ZN => n10075);
   U9546 : OAI22_X1 port map( A1 => n8795, A2 => n11689, B1 => n9243, B2 => 
                           n11685, ZN => n10083);
   U9547 : NAND4_X1 port map( A1 => n10084, A2 => n10085, A3 => n10086, A4 => 
                           n10087, ZN => n10082);
   U9548 : AOI221_X1 port map( B1 => n11626, B2 => n10867, C1 => n11622, C2 => 
                           n10739, A => n10091, ZN => n10084);
   U9549 : AOI221_X1 port map( B1 => n11696, B2 => n10065, C1 => n11693, C2 => 
                           Out2_23_port, A => n10066, ZN => n10058);
   U9550 : OAI22_X1 port map( A1 => n8794, A2 => n11689, B1 => n9242, B2 => 
                           n11685, ZN => n10066);
   U9551 : NAND4_X1 port map( A1 => n10067, A2 => n10068, A3 => n10069, A4 => 
                           n10070, ZN => n10065);
   U9552 : AOI221_X1 port map( B1 => n11626, B2 => n10868, C1 => n11622, C2 => 
                           n10740, A => n10074, ZN => n10067);
   U9553 : AOI221_X1 port map( B1 => n11696, B2 => n10048, C1 => n11693, C2 => 
                           Out2_24_port, A => n10049, ZN => n10041);
   U9554 : OAI22_X1 port map( A1 => n8793, A2 => n11690, B1 => n9241, B2 => 
                           n11686, ZN => n10049);
   U9555 : NAND4_X1 port map( A1 => n10050, A2 => n10051, A3 => n10052, A4 => 
                           n10053, ZN => n10048);
   U9556 : AOI221_X1 port map( B1 => n11627, B2 => n10869, C1 => n11623, C2 => 
                           n10741, A => n10057, ZN => n10050);
   U9557 : AOI221_X1 port map( B1 => n11696, B2 => n10031, C1 => n11694, C2 => 
                           Out2_25_port, A => n10032, ZN => n10024);
   U9558 : OAI22_X1 port map( A1 => n8792, A2 => n11690, B1 => n9240, B2 => 
                           n11686, ZN => n10032);
   U9559 : NAND4_X1 port map( A1 => n10033, A2 => n10034, A3 => n10035, A4 => 
                           n10036, ZN => n10031);
   U9560 : AOI221_X1 port map( B1 => n11627, B2 => n10870, C1 => n11623, C2 => 
                           n10742, A => n10040, ZN => n10033);
   U9561 : AOI221_X1 port map( B1 => n11696, B2 => n10014, C1 => n11694, C2 => 
                           Out2_26_port, A => n10015, ZN => n10007);
   U9562 : OAI22_X1 port map( A1 => n8791, A2 => n11690, B1 => n9239, B2 => 
                           n11686, ZN => n10015);
   U9563 : NAND4_X1 port map( A1 => n10016, A2 => n10017, A3 => n10018, A4 => 
                           n10019, ZN => n10014);
   U9564 : AOI221_X1 port map( B1 => n11627, B2 => n10871, C1 => n11623, C2 => 
                           n10743, A => n10023, ZN => n10016);
   U9565 : AOI221_X1 port map( B1 => n11696, B2 => n9997, C1 => n11694, C2 => 
                           Out2_27_port, A => n9998, ZN => n9990);
   U9566 : OAI22_X1 port map( A1 => n8790, A2 => n11690, B1 => n9238, B2 => 
                           n11686, ZN => n9998);
   U9567 : NAND4_X1 port map( A1 => n9999, A2 => n10000, A3 => n10001, A4 => 
                           n10002, ZN => n9997);
   U9568 : AOI221_X1 port map( B1 => n11627, B2 => n10872, C1 => n11623, C2 => 
                           n10744, A => n10006, ZN => n9999);
   U9569 : AOI221_X1 port map( B1 => n11696, B2 => n9980, C1 => n11694, C2 => 
                           Out2_28_port, A => n9981, ZN => n9973);
   U9570 : OAI22_X1 port map( A1 => n8789, A2 => n11690, B1 => n9237, B2 => 
                           n11686, ZN => n9981);
   U9571 : NAND4_X1 port map( A1 => n9982, A2 => n9983, A3 => n9984, A4 => 
                           n9985, ZN => n9980);
   U9572 : AOI221_X1 port map( B1 => n11627, B2 => n10873, C1 => n11623, C2 => 
                           n10745, A => n9989, ZN => n9982);
   U9573 : AOI221_X1 port map( B1 => n11696, B2 => n9963, C1 => n11694, C2 => 
                           Out2_29_port, A => n9964, ZN => n9956);
   U9574 : OAI22_X1 port map( A1 => n8788, A2 => n11690, B1 => n9236, B2 => 
                           n11686, ZN => n9964);
   U9575 : NAND4_X1 port map( A1 => n9965, A2 => n9966, A3 => n9967, A4 => 
                           n9968, ZN => n9963);
   U9576 : AOI221_X1 port map( B1 => n11627, B2 => n10874, C1 => n11623, C2 => 
                           n10746, A => n9972, ZN => n9965);
   U9577 : AOI221_X1 port map( B1 => n11696, B2 => n9946, C1 => n11694, C2 => 
                           Out2_30_port, A => n9947, ZN => n9939);
   U9578 : OAI22_X1 port map( A1 => n8787, A2 => n11690, B1 => n9235, B2 => 
                           n11686, ZN => n9947);
   U9579 : NAND4_X1 port map( A1 => n9948, A2 => n9949, A3 => n9950, A4 => 
                           n9951, ZN => n9946);
   U9580 : AOI221_X1 port map( B1 => n11627, B2 => n10875, C1 => n11623, C2 => 
                           n10747, A => n9955, ZN => n9948);
   U9581 : AOI221_X1 port map( B1 => n11696, B2 => n9908, C1 => n11694, C2 => 
                           Out2_31_port, A => n9910, ZN => n9888);
   U9582 : OAI22_X1 port map( A1 => n8786, A2 => n11690, B1 => n9234, B2 => 
                           n11686, ZN => n9910);
   U9583 : NAND4_X1 port map( A1 => n9913, A2 => n9914, A3 => n9915, A4 => 
                           n9916, ZN => n9908);
   U9584 : AOI221_X1 port map( B1 => n11627, B2 => n10876, C1 => n11623, C2 => 
                           n10748, A => n9936, ZN => n9913);
   U9585 : NAND4_X1 port map( A1 => n10449, A2 => n10450, A3 => n10451, A4 => 
                           n10452, ZN => n7214);
   U9586 : AOI221_X1 port map( B1 => n11716, B2 => n7398, C1 => n11712, C2 => 
                           n7558, A => n10462, ZN => n10450);
   U9587 : AOI221_X1 port map( B1 => n11732, B2 => n7590, C1 => n11728, C2 => 
                           n10909, A => n10459, ZN => n10451);
   U9588 : AOI221_X1 port map( B1 => n11748, B2 => n7494, C1 => n11744, C2 => 
                           n10941, A => n10453, ZN => n10452);
   U9589 : NAND4_X1 port map( A1 => n10432, A2 => n10433, A3 => n10434, A4 => 
                           n10435, ZN => n7215);
   U9590 : AOI221_X1 port map( B1 => n11716, B2 => n7399, C1 => n11712, C2 => 
                           n7559, A => n10438, ZN => n10433);
   U9591 : AOI221_X1 port map( B1 => n11732, B2 => n7591, C1 => n11728, C2 => 
                           n10910, A => n10437, ZN => n10434);
   U9592 : AOI221_X1 port map( B1 => n11748, B2 => n7495, C1 => n11744, C2 => 
                           n10942, A => n10436, ZN => n10435);
   U9593 : NAND4_X1 port map( A1 => n10415, A2 => n10416, A3 => n10417, A4 => 
                           n10418, ZN => n7216);
   U9594 : AOI221_X1 port map( B1 => n11716, B2 => n7400, C1 => n11712, C2 => 
                           n7560, A => n10421, ZN => n10416);
   U9595 : AOI221_X1 port map( B1 => n11732, B2 => n7592, C1 => n11728, C2 => 
                           n10911, A => n10420, ZN => n10417);
   U9596 : AOI221_X1 port map( B1 => n11748, B2 => n7496, C1 => n11744, C2 => 
                           n10943, A => n10419, ZN => n10418);
   U9597 : NAND4_X1 port map( A1 => n10398, A2 => n10399, A3 => n10400, A4 => 
                           n10401, ZN => n7217);
   U9598 : AOI221_X1 port map( B1 => n11716, B2 => n7401, C1 => n11712, C2 => 
                           n7561, A => n10404, ZN => n10399);
   U9599 : AOI221_X1 port map( B1 => n11732, B2 => n7593, C1 => n11728, C2 => 
                           n10912, A => n10403, ZN => n10400);
   U9600 : AOI221_X1 port map( B1 => n11748, B2 => n7497, C1 => n11744, C2 => 
                           n10944, A => n10402, ZN => n10401);
   U9601 : NAND4_X1 port map( A1 => n10381, A2 => n10382, A3 => n10383, A4 => 
                           n10384, ZN => n7218);
   U9602 : AOI221_X1 port map( B1 => n11716, B2 => n7402, C1 => n11712, C2 => 
                           n7562, A => n10387, ZN => n10382);
   U9603 : AOI221_X1 port map( B1 => n11732, B2 => n7594, C1 => n11728, C2 => 
                           n10913, A => n10386, ZN => n10383);
   U9604 : AOI221_X1 port map( B1 => n11748, B2 => n7498, C1 => n11744, C2 => 
                           n10945, A => n10385, ZN => n10384);
   U9605 : NAND4_X1 port map( A1 => n10364, A2 => n10365, A3 => n10366, A4 => 
                           n10367, ZN => n7219);
   U9606 : AOI221_X1 port map( B1 => n11716, B2 => n7403, C1 => n11712, C2 => 
                           n7563, A => n10370, ZN => n10365);
   U9607 : AOI221_X1 port map( B1 => n11732, B2 => n7595, C1 => n11728, C2 => 
                           n10914, A => n10369, ZN => n10366);
   U9608 : AOI221_X1 port map( B1 => n11748, B2 => n7499, C1 => n11744, C2 => 
                           n10946, A => n10368, ZN => n10367);
   U9609 : NAND4_X1 port map( A1 => n10347, A2 => n10348, A3 => n10349, A4 => 
                           n10350, ZN => n7220);
   U9610 : AOI221_X1 port map( B1 => n11716, B2 => n7404, C1 => n11712, C2 => 
                           n7564, A => n10353, ZN => n10348);
   U9611 : AOI221_X1 port map( B1 => n11732, B2 => n7596, C1 => n11728, C2 => 
                           n10915, A => n10352, ZN => n10349);
   U9612 : AOI221_X1 port map( B1 => n11748, B2 => n7500, C1 => n11744, C2 => 
                           n10947, A => n10351, ZN => n10350);
   U9613 : NAND4_X1 port map( A1 => n10330, A2 => n10331, A3 => n10332, A4 => 
                           n10333, ZN => n7221);
   U9614 : AOI221_X1 port map( B1 => n11716, B2 => n7405, C1 => n11712, C2 => 
                           n7565, A => n10336, ZN => n10331);
   U9615 : AOI221_X1 port map( B1 => n11732, B2 => n7597, C1 => n11728, C2 => 
                           n10916, A => n10335, ZN => n10332);
   U9616 : AOI221_X1 port map( B1 => n11748, B2 => n7501, C1 => n11744, C2 => 
                           n10948, A => n10334, ZN => n10333);
   U9617 : NAND4_X1 port map( A1 => n10313, A2 => n10314, A3 => n10315, A4 => 
                           n10316, ZN => n7222);
   U9618 : AOI221_X1 port map( B1 => n11716, B2 => n7397, C1 => n11712, C2 => 
                           n7557, A => n10319, ZN => n10314);
   U9619 : AOI221_X1 port map( B1 => n11732, B2 => n7589, C1 => n11728, C2 => 
                           n10917, A => n10318, ZN => n10315);
   U9620 : AOI221_X1 port map( B1 => n11748, B2 => n7493, C1 => n11744, C2 => 
                           n10949, A => n10317, ZN => n10316);
   U9621 : NAND4_X1 port map( A1 => n10296, A2 => n10297, A3 => n10298, A4 => 
                           n10299, ZN => n7223);
   U9622 : AOI221_X1 port map( B1 => n11716, B2 => n7374, C1 => n11712, C2 => 
                           n7534, A => n10302, ZN => n10297);
   U9623 : AOI221_X1 port map( B1 => n11732, B2 => n7566, C1 => n11728, C2 => 
                           n10918, A => n10301, ZN => n10298);
   U9624 : AOI221_X1 port map( B1 => n11748, B2 => n7470, C1 => n11744, C2 => 
                           n10950, A => n10300, ZN => n10299);
   U9625 : NAND4_X1 port map( A1 => n10279, A2 => n10280, A3 => n10281, A4 => 
                           n10282, ZN => n7224);
   U9626 : AOI221_X1 port map( B1 => n11716, B2 => n7375, C1 => n11712, C2 => 
                           n7535, A => n10285, ZN => n10280);
   U9627 : AOI221_X1 port map( B1 => n11732, B2 => n7567, C1 => n11728, C2 => 
                           n10919, A => n10284, ZN => n10281);
   U9628 : AOI221_X1 port map( B1 => n11748, B2 => n7471, C1 => n11744, C2 => 
                           n10951, A => n10283, ZN => n10282);
   U9629 : NAND4_X1 port map( A1 => n10262, A2 => n10263, A3 => n10264, A4 => 
                           n10265, ZN => n7225);
   U9630 : AOI221_X1 port map( B1 => n11716, B2 => n7376, C1 => n11712, C2 => 
                           n7536, A => n10268, ZN => n10263);
   U9631 : AOI221_X1 port map( B1 => n11732, B2 => n7568, C1 => n11728, C2 => 
                           n10920, A => n10267, ZN => n10264);
   U9632 : AOI221_X1 port map( B1 => n11748, B2 => n7472, C1 => n11744, C2 => 
                           n10952, A => n10266, ZN => n10265);
   U9633 : NAND4_X1 port map( A1 => n10245, A2 => n10246, A3 => n10247, A4 => 
                           n10248, ZN => n7226);
   U9634 : AOI221_X1 port map( B1 => n11717, B2 => n7377, C1 => n11713, C2 => 
                           n7537, A => n10251, ZN => n10246);
   U9635 : AOI221_X1 port map( B1 => n11733, B2 => n7569, C1 => n11729, C2 => 
                           n10921, A => n10250, ZN => n10247);
   U9636 : AOI221_X1 port map( B1 => n11749, B2 => n7473, C1 => n11745, C2 => 
                           n10953, A => n10249, ZN => n10248);
   U9637 : NAND4_X1 port map( A1 => n10228, A2 => n10229, A3 => n10230, A4 => 
                           n10231, ZN => n7227);
   U9638 : AOI221_X1 port map( B1 => n11717, B2 => n7378, C1 => n11713, C2 => 
                           n7538, A => n10234, ZN => n10229);
   U9639 : AOI221_X1 port map( B1 => n11733, B2 => n7570, C1 => n11729, C2 => 
                           n10922, A => n10233, ZN => n10230);
   U9640 : AOI221_X1 port map( B1 => n11749, B2 => n7474, C1 => n11745, C2 => 
                           n10954, A => n10232, ZN => n10231);
   U9641 : NAND4_X1 port map( A1 => n10211, A2 => n10212, A3 => n10213, A4 => 
                           n10214, ZN => n7228);
   U9642 : AOI221_X1 port map( B1 => n11717, B2 => n7379, C1 => n11713, C2 => 
                           n7539, A => n10217, ZN => n10212);
   U9643 : AOI221_X1 port map( B1 => n11733, B2 => n7571, C1 => n11729, C2 => 
                           n10923, A => n10216, ZN => n10213);
   U9644 : AOI221_X1 port map( B1 => n11749, B2 => n7475, C1 => n11745, C2 => 
                           n10955, A => n10215, ZN => n10214);
   U9645 : NAND4_X1 port map( A1 => n10194, A2 => n10195, A3 => n10196, A4 => 
                           n10197, ZN => n7229);
   U9646 : AOI221_X1 port map( B1 => n11717, B2 => n7380, C1 => n11713, C2 => 
                           n7540, A => n10200, ZN => n10195);
   U9647 : AOI221_X1 port map( B1 => n11733, B2 => n7572, C1 => n11729, C2 => 
                           n10924, A => n10199, ZN => n10196);
   U9648 : AOI221_X1 port map( B1 => n11749, B2 => n7476, C1 => n11745, C2 => 
                           n10956, A => n10198, ZN => n10197);
   U9649 : NAND4_X1 port map( A1 => n10177, A2 => n10178, A3 => n10179, A4 => 
                           n10180, ZN => n7230);
   U9650 : AOI221_X1 port map( B1 => n11717, B2 => n7381, C1 => n11713, C2 => 
                           n7541, A => n10183, ZN => n10178);
   U9651 : AOI221_X1 port map( B1 => n11733, B2 => n7573, C1 => n11729, C2 => 
                           n10925, A => n10182, ZN => n10179);
   U9652 : AOI221_X1 port map( B1 => n11749, B2 => n7477, C1 => n11745, C2 => 
                           n10957, A => n10181, ZN => n10180);
   U9653 : NAND4_X1 port map( A1 => n10160, A2 => n10161, A3 => n10162, A4 => 
                           n10163, ZN => n7231);
   U9654 : AOI221_X1 port map( B1 => n11717, B2 => n7382, C1 => n11713, C2 => 
                           n7542, A => n10166, ZN => n10161);
   U9655 : AOI221_X1 port map( B1 => n11733, B2 => n7574, C1 => n11729, C2 => 
                           n10926, A => n10165, ZN => n10162);
   U9656 : AOI221_X1 port map( B1 => n11749, B2 => n7478, C1 => n11745, C2 => 
                           n10958, A => n10164, ZN => n10163);
   U9657 : NAND4_X1 port map( A1 => n10143, A2 => n10144, A3 => n10145, A4 => 
                           n10146, ZN => n7232);
   U9658 : AOI221_X1 port map( B1 => n11717, B2 => n7383, C1 => n11713, C2 => 
                           n7543, A => n10149, ZN => n10144);
   U9659 : AOI221_X1 port map( B1 => n11733, B2 => n7575, C1 => n11729, C2 => 
                           n10927, A => n10148, ZN => n10145);
   U9660 : AOI221_X1 port map( B1 => n11749, B2 => n7479, C1 => n11745, C2 => 
                           n10959, A => n10147, ZN => n10146);
   U9661 : NAND4_X1 port map( A1 => n10126, A2 => n10127, A3 => n10128, A4 => 
                           n10129, ZN => n7233);
   U9662 : AOI221_X1 port map( B1 => n11717, B2 => n7384, C1 => n11713, C2 => 
                           n7544, A => n10132, ZN => n10127);
   U9663 : AOI221_X1 port map( B1 => n11733, B2 => n7576, C1 => n11729, C2 => 
                           n10928, A => n10131, ZN => n10128);
   U9664 : AOI221_X1 port map( B1 => n11749, B2 => n7480, C1 => n11745, C2 => 
                           n10960, A => n10130, ZN => n10129);
   U9665 : NAND4_X1 port map( A1 => n10109, A2 => n10110, A3 => n10111, A4 => 
                           n10112, ZN => n7234);
   U9666 : AOI221_X1 port map( B1 => n11717, B2 => n7385, C1 => n11713, C2 => 
                           n7545, A => n10115, ZN => n10110);
   U9667 : AOI221_X1 port map( B1 => n11733, B2 => n7577, C1 => n11729, C2 => 
                           n10929, A => n10114, ZN => n10111);
   U9668 : AOI221_X1 port map( B1 => n11749, B2 => n7481, C1 => n11745, C2 => 
                           n10961, A => n10113, ZN => n10112);
   U9669 : NAND4_X1 port map( A1 => n10092, A2 => n10093, A3 => n10094, A4 => 
                           n10095, ZN => n7235);
   U9670 : AOI221_X1 port map( B1 => n11717, B2 => n7386, C1 => n11713, C2 => 
                           n7546, A => n10098, ZN => n10093);
   U9671 : AOI221_X1 port map( B1 => n11733, B2 => n7578, C1 => n11729, C2 => 
                           n10930, A => n10097, ZN => n10094);
   U9672 : AOI221_X1 port map( B1 => n11749, B2 => n7482, C1 => n11745, C2 => 
                           n10962, A => n10096, ZN => n10095);
   U9673 : NAND4_X1 port map( A1 => n10075, A2 => n10076, A3 => n10077, A4 => 
                           n10078, ZN => n7236);
   U9674 : AOI221_X1 port map( B1 => n11717, B2 => n7387, C1 => n11713, C2 => 
                           n7547, A => n10081, ZN => n10076);
   U9675 : AOI221_X1 port map( B1 => n11733, B2 => n7579, C1 => n11729, C2 => 
                           n10931, A => n10080, ZN => n10077);
   U9676 : AOI221_X1 port map( B1 => n11749, B2 => n7483, C1 => n11745, C2 => 
                           n10963, A => n10079, ZN => n10078);
   U9677 : NAND4_X1 port map( A1 => n10058, A2 => n10059, A3 => n10060, A4 => 
                           n10061, ZN => n7237);
   U9678 : AOI221_X1 port map( B1 => n11717, B2 => n7388, C1 => n11713, C2 => 
                           n7548, A => n10064, ZN => n10059);
   U9679 : AOI221_X1 port map( B1 => n11733, B2 => n7580, C1 => n11729, C2 => 
                           n10932, A => n10063, ZN => n10060);
   U9680 : AOI221_X1 port map( B1 => n11749, B2 => n7484, C1 => n11745, C2 => 
                           n10964, A => n10062, ZN => n10061);
   U9681 : NAND4_X1 port map( A1 => n10041, A2 => n10042, A3 => n10043, A4 => 
                           n10044, ZN => n7238);
   U9682 : AOI221_X1 port map( B1 => n11718, B2 => n7389, C1 => n11714, C2 => 
                           n7549, A => n10047, ZN => n10042);
   U9683 : AOI221_X1 port map( B1 => n11734, B2 => n7581, C1 => n11730, C2 => 
                           n10933, A => n10046, ZN => n10043);
   U9684 : AOI221_X1 port map( B1 => n11750, B2 => n7485, C1 => n11746, C2 => 
                           n10965, A => n10045, ZN => n10044);
   U9685 : NAND4_X1 port map( A1 => n10024, A2 => n10025, A3 => n10026, A4 => 
                           n10027, ZN => n7239);
   U9686 : AOI221_X1 port map( B1 => n11718, B2 => n7390, C1 => n11714, C2 => 
                           n7550, A => n10030, ZN => n10025);
   U9687 : AOI221_X1 port map( B1 => n11734, B2 => n7582, C1 => n11730, C2 => 
                           n10934, A => n10029, ZN => n10026);
   U9688 : AOI221_X1 port map( B1 => n11750, B2 => n7486, C1 => n11746, C2 => 
                           n10966, A => n10028, ZN => n10027);
   U9689 : NAND4_X1 port map( A1 => n10007, A2 => n10008, A3 => n10009, A4 => 
                           n10010, ZN => n7240);
   U9690 : AOI221_X1 port map( B1 => n11718, B2 => n7391, C1 => n11714, C2 => 
                           n7551, A => n10013, ZN => n10008);
   U9691 : AOI221_X1 port map( B1 => n11734, B2 => n7583, C1 => n11730, C2 => 
                           n10935, A => n10012, ZN => n10009);
   U9692 : AOI221_X1 port map( B1 => n11750, B2 => n7487, C1 => n11746, C2 => 
                           n10967, A => n10011, ZN => n10010);
   U9693 : NAND4_X1 port map( A1 => n9990, A2 => n9991, A3 => n9992, A4 => 
                           n9993, ZN => n7241);
   U9694 : AOI221_X1 port map( B1 => n11718, B2 => n7392, C1 => n11714, C2 => 
                           n7552, A => n9996, ZN => n9991);
   U9695 : AOI221_X1 port map( B1 => n11734, B2 => n7584, C1 => n11730, C2 => 
                           n10936, A => n9995, ZN => n9992);
   U9696 : AOI221_X1 port map( B1 => n11750, B2 => n7488, C1 => n11746, C2 => 
                           n10968, A => n9994, ZN => n9993);
   U9697 : NAND4_X1 port map( A1 => n9973, A2 => n9974, A3 => n9975, A4 => 
                           n9976, ZN => n7242);
   U9698 : AOI221_X1 port map( B1 => n11718, B2 => n7393, C1 => n11714, C2 => 
                           n7553, A => n9979, ZN => n9974);
   U9699 : AOI221_X1 port map( B1 => n11734, B2 => n7585, C1 => n11730, C2 => 
                           n10937, A => n9978, ZN => n9975);
   U9700 : AOI221_X1 port map( B1 => n11750, B2 => n7489, C1 => n11746, C2 => 
                           n10969, A => n9977, ZN => n9976);
   U9701 : NAND4_X1 port map( A1 => n9956, A2 => n9957, A3 => n9958, A4 => 
                           n9959, ZN => n7243);
   U9702 : AOI221_X1 port map( B1 => n11718, B2 => n7394, C1 => n11714, C2 => 
                           n7554, A => n9962, ZN => n9957);
   U9703 : AOI221_X1 port map( B1 => n11734, B2 => n7586, C1 => n11730, C2 => 
                           n10938, A => n9961, ZN => n9958);
   U9704 : AOI221_X1 port map( B1 => n11750, B2 => n7490, C1 => n11746, C2 => 
                           n10970, A => n9960, ZN => n9959);
   U9705 : NAND4_X1 port map( A1 => n9939, A2 => n9940, A3 => n9941, A4 => 
                           n9942, ZN => n7244);
   U9706 : AOI221_X1 port map( B1 => n11718, B2 => n7395, C1 => n11714, C2 => 
                           n7555, A => n9945, ZN => n9940);
   U9707 : AOI221_X1 port map( B1 => n11734, B2 => n7587, C1 => n11730, C2 => 
                           n10939, A => n9944, ZN => n9941);
   U9708 : AOI221_X1 port map( B1 => n11750, B2 => n7491, C1 => n11746, C2 => 
                           n10971, A => n9943, ZN => n9942);
   U9709 : NAND4_X1 port map( A1 => n9888, A2 => n9889, A3 => n9890, A4 => 
                           n9891, ZN => n7245);
   U9710 : AOI221_X1 port map( B1 => n11718, B2 => n7396, C1 => n11714, C2 => 
                           n7556, A => n9904, ZN => n9889);
   U9711 : AOI221_X1 port map( B1 => n11734, B2 => n7588, C1 => n11730, C2 => 
                           n10940, A => n9899, ZN => n9890);
   U9712 : AOI221_X1 port map( B1 => n11750, B2 => n7492, C1 => n11746, C2 => 
                           n10972, A => n9894, ZN => n9891);
   U9713 : AOI221_X1 port map( B1 => n11133, B2 => n11784, C1 => n11005, C2 => 
                           n11780, A => n9886, ZN => n9878);
   U9714 : OAI222_X1 port map( A1 => n11776, A2 => n8369, B1 => n11772, B2 => 
                           n8689, C1 => n11768, C2 => n8625, ZN => n9886);
   U9715 : AOI221_X1 port map( B1 => n11134, B2 => n11784, C1 => n11006, C2 => 
                           n11780, A => n9857, ZN => n9852);
   U9716 : OAI222_X1 port map( A1 => n11776, A2 => n8368, B1 => n11772, B2 => 
                           n8688, C1 => n11768, C2 => n8624, ZN => n9857);
   U9717 : AOI221_X1 port map( B1 => n11135, B2 => n11784, C1 => n11007, C2 => 
                           n11780, A => n9840, ZN => n9835);
   U9718 : OAI222_X1 port map( A1 => n11776, A2 => n8367, B1 => n11772, B2 => 
                           n8687, C1 => n11768, C2 => n8623, ZN => n9840);
   U9719 : AOI221_X1 port map( B1 => n11136, B2 => n11784, C1 => n11008, C2 => 
                           n11780, A => n9823, ZN => n9818);
   U9720 : OAI222_X1 port map( A1 => n11776, A2 => n8366, B1 => n11772, B2 => 
                           n8686, C1 => n11768, C2 => n8622, ZN => n9823);
   U9721 : AOI221_X1 port map( B1 => n11137, B2 => n11784, C1 => n11009, C2 => 
                           n11780, A => n9806, ZN => n9801);
   U9722 : OAI222_X1 port map( A1 => n11776, A2 => n8365, B1 => n11772, B2 => 
                           n8685, C1 => n11768, C2 => n8621, ZN => n9806);
   U9723 : AOI221_X1 port map( B1 => n11138, B2 => n11784, C1 => n11010, C2 => 
                           n11780, A => n9789, ZN => n9784);
   U9724 : OAI222_X1 port map( A1 => n11776, A2 => n8364, B1 => n11772, B2 => 
                           n8684, C1 => n11768, C2 => n8620, ZN => n9789);
   U9725 : AOI221_X1 port map( B1 => n11139, B2 => n11784, C1 => n11011, C2 => 
                           n11780, A => n9772, ZN => n9767);
   U9726 : OAI222_X1 port map( A1 => n11776, A2 => n8363, B1 => n11772, B2 => 
                           n8683, C1 => n11768, C2 => n8619, ZN => n9772);
   U9727 : AOI221_X1 port map( B1 => n11140, B2 => n11784, C1 => n11012, C2 => 
                           n11780, A => n9755, ZN => n9750);
   U9728 : OAI222_X1 port map( A1 => n11776, A2 => n8362, B1 => n11772, B2 => 
                           n8682, C1 => n11768, C2 => n8618, ZN => n9755);
   U9729 : AOI221_X1 port map( B1 => n11141, B2 => n11784, C1 => n11013, C2 => 
                           n11780, A => n9738, ZN => n9733);
   U9730 : OAI222_X1 port map( A1 => n11776, A2 => n8361, B1 => n11772, B2 => 
                           n8681, C1 => n11768, C2 => n8617, ZN => n9738);
   U9731 : AOI221_X1 port map( B1 => n11142, B2 => n11784, C1 => n11014, C2 => 
                           n11780, A => n9721, ZN => n9716);
   U9732 : OAI222_X1 port map( A1 => n11776, A2 => n8360, B1 => n11772, B2 => 
                           n8680, C1 => n11768, C2 => n8616, ZN => n9721);
   U9733 : AOI221_X1 port map( B1 => n11143, B2 => n11784, C1 => n11015, C2 => 
                           n11780, A => n9704, ZN => n9699);
   U9734 : OAI222_X1 port map( A1 => n11776, A2 => n8359, B1 => n11772, B2 => 
                           n8679, C1 => n11768, C2 => n8615, ZN => n9704);
   U9735 : AOI221_X1 port map( B1 => n11144, B2 => n11784, C1 => n11016, C2 => 
                           n11780, A => n9687, ZN => n9682);
   U9736 : OAI222_X1 port map( A1 => n11776, A2 => n8358, B1 => n11772, B2 => 
                           n8678, C1 => n11768, C2 => n8614, ZN => n9687);
   U9737 : AOI221_X1 port map( B1 => n11145, B2 => n11785, C1 => n11017, C2 => 
                           n11781, A => n9670, ZN => n9665);
   U9738 : OAI222_X1 port map( A1 => n11777, A2 => n8357, B1 => n11773, B2 => 
                           n8677, C1 => n11769, C2 => n8613, ZN => n9670);
   U9739 : AOI221_X1 port map( B1 => n11146, B2 => n11785, C1 => n11018, C2 => 
                           n11781, A => n9653, ZN => n9648);
   U9740 : OAI222_X1 port map( A1 => n11777, A2 => n8356, B1 => n11773, B2 => 
                           n8676, C1 => n11769, C2 => n8612, ZN => n9653);
   U9741 : AOI221_X1 port map( B1 => n11147, B2 => n11785, C1 => n11019, C2 => 
                           n11781, A => n9636, ZN => n9631);
   U9742 : OAI222_X1 port map( A1 => n11777, A2 => n8355, B1 => n11773, B2 => 
                           n8675, C1 => n11769, C2 => n8611, ZN => n9636);
   U9743 : AOI221_X1 port map( B1 => n11148, B2 => n11785, C1 => n11020, C2 => 
                           n11781, A => n9619, ZN => n9614);
   U9744 : OAI222_X1 port map( A1 => n11777, A2 => n8354, B1 => n11773, B2 => 
                           n8674, C1 => n11769, C2 => n8610, ZN => n9619);
   U9745 : AOI221_X1 port map( B1 => n11149, B2 => n11785, C1 => n11021, C2 => 
                           n11781, A => n9602, ZN => n9597);
   U9746 : OAI222_X1 port map( A1 => n11777, A2 => n8353, B1 => n11773, B2 => 
                           n8673, C1 => n11769, C2 => n8609, ZN => n9602);
   U9747 : AOI221_X1 port map( B1 => n11150, B2 => n11785, C1 => n11022, C2 => 
                           n11781, A => n9585, ZN => n9580);
   U9748 : OAI222_X1 port map( A1 => n11777, A2 => n8352, B1 => n11773, B2 => 
                           n8672, C1 => n11769, C2 => n8608, ZN => n9585);
   U9749 : AOI221_X1 port map( B1 => n11151, B2 => n11785, C1 => n11023, C2 => 
                           n11781, A => n9568, ZN => n9563);
   U9750 : OAI222_X1 port map( A1 => n11777, A2 => n8351, B1 => n11773, B2 => 
                           n8671, C1 => n11769, C2 => n8607, ZN => n9568);
   U9751 : AOI221_X1 port map( B1 => n11152, B2 => n11785, C1 => n11024, C2 => 
                           n11781, A => n9551, ZN => n9546);
   U9752 : OAI222_X1 port map( A1 => n11777, A2 => n8350, B1 => n11773, B2 => 
                           n8670, C1 => n11769, C2 => n8606, ZN => n9551);
   U9753 : AOI221_X1 port map( B1 => n11153, B2 => n11785, C1 => n11025, C2 => 
                           n11781, A => n9534, ZN => n9529);
   U9754 : OAI222_X1 port map( A1 => n11777, A2 => n8349, B1 => n11773, B2 => 
                           n8669, C1 => n11769, C2 => n8605, ZN => n9534);
   U9755 : AOI221_X1 port map( B1 => n11154, B2 => n11785, C1 => n11026, C2 => 
                           n11781, A => n9517, ZN => n9512);
   U9756 : OAI222_X1 port map( A1 => n11777, A2 => n8348, B1 => n11773, B2 => 
                           n8668, C1 => n11769, C2 => n8604, ZN => n9517);
   U9757 : AOI221_X1 port map( B1 => n11155, B2 => n11785, C1 => n11027, C2 => 
                           n11781, A => n9500, ZN => n9495);
   U9758 : OAI222_X1 port map( A1 => n11777, A2 => n8347, B1 => n11773, B2 => 
                           n8667, C1 => n11769, C2 => n8603, ZN => n9500);
   U9759 : AOI221_X1 port map( B1 => n11156, B2 => n11785, C1 => n11028, C2 => 
                           n11781, A => n9483, ZN => n9478);
   U9760 : OAI222_X1 port map( A1 => n11777, A2 => n8346, B1 => n11773, B2 => 
                           n8666, C1 => n11769, C2 => n8602, ZN => n9483);
   U9761 : AOI221_X1 port map( B1 => n11157, B2 => n11786, C1 => n11029, C2 => 
                           n11782, A => n9466, ZN => n9461);
   U9762 : OAI222_X1 port map( A1 => n11778, A2 => n8345, B1 => n11774, B2 => 
                           n8665, C1 => n11770, C2 => n8601, ZN => n9466);
   U9763 : AOI221_X1 port map( B1 => n11158, B2 => n11786, C1 => n11030, C2 => 
                           n11782, A => n9449, ZN => n9444);
   U9764 : OAI222_X1 port map( A1 => n11778, A2 => n8344, B1 => n11774, B2 => 
                           n8664, C1 => n11770, C2 => n8600, ZN => n9449);
   U9765 : AOI221_X1 port map( B1 => n11159, B2 => n11786, C1 => n11031, C2 => 
                           n11782, A => n9432, ZN => n9427);
   U9766 : OAI222_X1 port map( A1 => n11778, A2 => n8343, B1 => n11774, B2 => 
                           n8663, C1 => n11770, C2 => n8599, ZN => n9432);
   U9767 : AOI221_X1 port map( B1 => n11160, B2 => n11786, C1 => n11032, C2 => 
                           n11782, A => n9415, ZN => n9410);
   U9768 : OAI222_X1 port map( A1 => n11778, A2 => n8342, B1 => n11774, B2 => 
                           n8662, C1 => n11770, C2 => n8598, ZN => n9415);
   U9769 : AOI221_X1 port map( B1 => n11161, B2 => n11786, C1 => n11033, C2 => 
                           n11782, A => n9398, ZN => n9393);
   U9770 : OAI222_X1 port map( A1 => n11778, A2 => n8341, B1 => n11774, B2 => 
                           n8661, C1 => n11770, C2 => n8597, ZN => n9398);
   U9771 : AOI221_X1 port map( B1 => n11162, B2 => n11786, C1 => n11034, C2 => 
                           n11782, A => n9381, ZN => n9376);
   U9772 : OAI222_X1 port map( A1 => n11778, A2 => n8340, B1 => n11774, B2 => 
                           n8660, C1 => n11770, C2 => n8596, ZN => n9381);
   U9773 : AOI221_X1 port map( B1 => n11163, B2 => n11786, C1 => n11035, C2 => 
                           n11782, A => n9364, ZN => n9359);
   U9774 : OAI222_X1 port map( A1 => n11778, A2 => n8339, B1 => n11774, B2 => 
                           n8659, C1 => n11770, C2 => n8595, ZN => n9364);
   U9775 : AOI221_X1 port map( B1 => n11164, B2 => n11786, C1 => n11036, C2 => 
                           n11782, A => n9340, ZN => n9324);
   U9776 : OAI222_X1 port map( A1 => n11778, A2 => n8338, B1 => n11774, B2 => 
                           n8658, C1 => n11770, C2 => n8594, ZN => n9340);
   U9777 : AOI221_X1 port map( B1 => n11647, B2 => n11157, C1 => n11643, C2 => 
                           n11029, A => n10056, ZN => n10051);
   U9778 : OAI222_X1 port map( A1 => n8345, A2 => n11639, B1 => n8665, B2 => 
                           n11635, C1 => n8601, C2 => n11631, ZN => n10056);
   U9779 : AOI221_X1 port map( B1 => n11647, B2 => n11158, C1 => n11643, C2 => 
                           n11030, A => n10039, ZN => n10034);
   U9780 : OAI222_X1 port map( A1 => n8344, A2 => n11639, B1 => n8664, B2 => 
                           n11635, C1 => n8600, C2 => n11631, ZN => n10039);
   U9781 : AOI221_X1 port map( B1 => n11647, B2 => n11159, C1 => n11643, C2 => 
                           n11031, A => n10022, ZN => n10017);
   U9782 : OAI222_X1 port map( A1 => n8343, A2 => n11639, B1 => n8663, B2 => 
                           n11635, C1 => n8599, C2 => n11631, ZN => n10022);
   U9783 : AOI221_X1 port map( B1 => n11647, B2 => n11160, C1 => n11643, C2 => 
                           n11032, A => n10005, ZN => n10000);
   U9784 : OAI222_X1 port map( A1 => n8342, A2 => n11639, B1 => n8662, B2 => 
                           n11635, C1 => n8598, C2 => n11631, ZN => n10005);
   U9785 : AOI221_X1 port map( B1 => n11647, B2 => n11161, C1 => n11643, C2 => 
                           n11033, A => n9988, ZN => n9983);
   U9786 : OAI222_X1 port map( A1 => n8341, A2 => n11639, B1 => n8661, B2 => 
                           n11635, C1 => n8597, C2 => n11631, ZN => n9988);
   U9787 : AOI221_X1 port map( B1 => n11647, B2 => n11162, C1 => n11643, C2 => 
                           n11034, A => n9971, ZN => n9966);
   U9788 : OAI222_X1 port map( A1 => n8340, A2 => n11639, B1 => n8660, B2 => 
                           n11635, C1 => n8596, C2 => n11631, ZN => n9971);
   U9789 : AOI221_X1 port map( B1 => n11647, B2 => n11163, C1 => n11643, C2 => 
                           n11035, A => n9954, ZN => n9949);
   U9790 : OAI222_X1 port map( A1 => n8339, A2 => n11639, B1 => n8659, B2 => 
                           n11635, C1 => n8595, C2 => n11631, ZN => n9954);
   U9791 : AOI221_X1 port map( B1 => n11647, B2 => n11164, C1 => n11643, C2 => 
                           n11036, A => n9930, ZN => n9914);
   U9792 : OAI222_X1 port map( A1 => n8338, A2 => n11639, B1 => n8658, B2 => 
                           n11635, C1 => n8594, C2 => n11631, ZN => n9930);
   U9793 : AOI221_X1 port map( B1 => n11645, B2 => n11133, C1 => n11641, C2 => 
                           n11005, A => n10476, ZN => n10468);
   U9794 : OAI222_X1 port map( A1 => n8369, A2 => n11637, B1 => n8689, B2 => 
                           n11633, C1 => n8625, C2 => n11629, ZN => n10476);
   U9795 : AOI221_X1 port map( B1 => n11645, B2 => n11134, C1 => n11641, C2 => 
                           n11006, A => n10447, ZN => n10442);
   U9796 : OAI222_X1 port map( A1 => n8368, A2 => n11637, B1 => n8688, B2 => 
                           n11633, C1 => n8624, C2 => n11629, ZN => n10447);
   U9797 : AOI221_X1 port map( B1 => n11645, B2 => n11135, C1 => n11641, C2 => 
                           n11007, A => n10430, ZN => n10425);
   U9798 : OAI222_X1 port map( A1 => n8367, A2 => n11637, B1 => n8687, B2 => 
                           n11633, C1 => n8623, C2 => n11629, ZN => n10430);
   U9799 : AOI221_X1 port map( B1 => n11645, B2 => n11136, C1 => n11641, C2 => 
                           n11008, A => n10413, ZN => n10408);
   U9800 : OAI222_X1 port map( A1 => n8366, A2 => n11637, B1 => n8686, B2 => 
                           n11633, C1 => n8622, C2 => n11629, ZN => n10413);
   U9801 : AOI221_X1 port map( B1 => n11645, B2 => n11137, C1 => n11641, C2 => 
                           n11009, A => n10396, ZN => n10391);
   U9802 : OAI222_X1 port map( A1 => n8365, A2 => n11637, B1 => n8685, B2 => 
                           n11633, C1 => n8621, C2 => n11629, ZN => n10396);
   U9803 : AOI221_X1 port map( B1 => n11645, B2 => n11138, C1 => n11641, C2 => 
                           n11010, A => n10379, ZN => n10374);
   U9804 : OAI222_X1 port map( A1 => n8364, A2 => n11637, B1 => n8684, B2 => 
                           n11633, C1 => n8620, C2 => n11629, ZN => n10379);
   U9805 : AOI221_X1 port map( B1 => n11645, B2 => n11139, C1 => n11641, C2 => 
                           n11011, A => n10362, ZN => n10357);
   U9806 : OAI222_X1 port map( A1 => n8363, A2 => n11637, B1 => n8683, B2 => 
                           n11633, C1 => n8619, C2 => n11629, ZN => n10362);
   U9807 : AOI221_X1 port map( B1 => n11645, B2 => n11140, C1 => n11641, C2 => 
                           n11012, A => n10345, ZN => n10340);
   U9808 : OAI222_X1 port map( A1 => n8362, A2 => n11637, B1 => n8682, B2 => 
                           n11633, C1 => n8618, C2 => n11629, ZN => n10345);
   U9809 : AOI221_X1 port map( B1 => n11645, B2 => n11141, C1 => n11641, C2 => 
                           n11013, A => n10328, ZN => n10323);
   U9810 : OAI222_X1 port map( A1 => n8361, A2 => n11637, B1 => n8681, B2 => 
                           n11633, C1 => n8617, C2 => n11629, ZN => n10328);
   U9811 : AOI221_X1 port map( B1 => n11645, B2 => n11142, C1 => n11641, C2 => 
                           n11014, A => n10311, ZN => n10306);
   U9812 : OAI222_X1 port map( A1 => n8360, A2 => n11637, B1 => n8680, B2 => 
                           n11633, C1 => n8616, C2 => n11629, ZN => n10311);
   U9813 : AOI221_X1 port map( B1 => n11645, B2 => n11143, C1 => n11641, C2 => 
                           n11015, A => n10294, ZN => n10289);
   U9814 : OAI222_X1 port map( A1 => n8359, A2 => n11637, B1 => n8679, B2 => 
                           n11633, C1 => n8615, C2 => n11629, ZN => n10294);
   U9815 : AOI221_X1 port map( B1 => n11645, B2 => n11144, C1 => n11641, C2 => 
                           n11016, A => n10277, ZN => n10272);
   U9816 : OAI222_X1 port map( A1 => n8358, A2 => n11637, B1 => n8678, B2 => 
                           n11633, C1 => n8614, C2 => n11629, ZN => n10277);
   U9817 : AOI221_X1 port map( B1 => n11646, B2 => n11145, C1 => n11642, C2 => 
                           n11017, A => n10260, ZN => n10255);
   U9818 : OAI222_X1 port map( A1 => n8357, A2 => n11638, B1 => n8677, B2 => 
                           n11634, C1 => n8613, C2 => n11630, ZN => n10260);
   U9819 : AOI221_X1 port map( B1 => n11646, B2 => n11146, C1 => n11642, C2 => 
                           n11018, A => n10243, ZN => n10238);
   U9820 : OAI222_X1 port map( A1 => n8356, A2 => n11638, B1 => n8676, B2 => 
                           n11634, C1 => n8612, C2 => n11630, ZN => n10243);
   U9821 : AOI221_X1 port map( B1 => n11646, B2 => n11147, C1 => n11642, C2 => 
                           n11019, A => n10226, ZN => n10221);
   U9822 : OAI222_X1 port map( A1 => n8355, A2 => n11638, B1 => n8675, B2 => 
                           n11634, C1 => n8611, C2 => n11630, ZN => n10226);
   U9823 : AOI221_X1 port map( B1 => n11646, B2 => n11148, C1 => n11642, C2 => 
                           n11020, A => n10209, ZN => n10204);
   U9824 : OAI222_X1 port map( A1 => n8354, A2 => n11638, B1 => n8674, B2 => 
                           n11634, C1 => n8610, C2 => n11630, ZN => n10209);
   U9825 : AOI221_X1 port map( B1 => n11646, B2 => n11149, C1 => n11642, C2 => 
                           n11021, A => n10192, ZN => n10187);
   U9826 : OAI222_X1 port map( A1 => n8353, A2 => n11638, B1 => n8673, B2 => 
                           n11634, C1 => n8609, C2 => n11630, ZN => n10192);
   U9827 : AOI221_X1 port map( B1 => n11646, B2 => n11150, C1 => n11642, C2 => 
                           n11022, A => n10175, ZN => n10170);
   U9828 : OAI222_X1 port map( A1 => n8352, A2 => n11638, B1 => n8672, B2 => 
                           n11634, C1 => n8608, C2 => n11630, ZN => n10175);
   U9829 : AOI221_X1 port map( B1 => n11646, B2 => n11151, C1 => n11642, C2 => 
                           n11023, A => n10158, ZN => n10153);
   U9830 : OAI222_X1 port map( A1 => n8351, A2 => n11638, B1 => n8671, B2 => 
                           n11634, C1 => n8607, C2 => n11630, ZN => n10158);
   U9831 : AOI221_X1 port map( B1 => n11646, B2 => n11152, C1 => n11642, C2 => 
                           n11024, A => n10141, ZN => n10136);
   U9832 : OAI222_X1 port map( A1 => n8350, A2 => n11638, B1 => n8670, B2 => 
                           n11634, C1 => n8606, C2 => n11630, ZN => n10141);
   U9833 : AOI221_X1 port map( B1 => n11646, B2 => n11153, C1 => n11642, C2 => 
                           n11025, A => n10124, ZN => n10119);
   U9834 : OAI222_X1 port map( A1 => n8349, A2 => n11638, B1 => n8669, B2 => 
                           n11634, C1 => n8605, C2 => n11630, ZN => n10124);
   U9835 : AOI221_X1 port map( B1 => n11646, B2 => n11154, C1 => n11642, C2 => 
                           n11026, A => n10107, ZN => n10102);
   U9836 : OAI222_X1 port map( A1 => n8348, A2 => n11638, B1 => n8668, B2 => 
                           n11634, C1 => n8604, C2 => n11630, ZN => n10107);
   U9837 : AOI221_X1 port map( B1 => n11646, B2 => n11155, C1 => n11642, C2 => 
                           n11027, A => n10090, ZN => n10085);
   U9838 : OAI222_X1 port map( A1 => n8347, A2 => n11638, B1 => n8667, B2 => 
                           n11634, C1 => n8603, C2 => n11630, ZN => n10090);
   U9839 : AOI221_X1 port map( B1 => n11646, B2 => n11156, C1 => n11642, C2 => 
                           n11028, A => n10073, ZN => n10068);
   U9840 : OAI222_X1 port map( A1 => n8346, A2 => n11638, B1 => n8666, B2 => 
                           n11634, C1 => n8602, C2 => n11630, ZN => n10073);
   U9841 : AOI221_X1 port map( B1 => n10973, B2 => n11800, C1 => n11165, C2 => 
                           n11796, A => n9885, ZN => n9879);
   U9842 : OAI22_X1 port map( A1 => n11792, A2 => n8433, B1 => n11788, B2 => 
                           n8657, ZN => n9885);
   U9843 : AOI221_X1 port map( B1 => n10974, B2 => n11800, C1 => n11166, C2 => 
                           n11796, A => n9856, ZN => n9853);
   U9844 : OAI22_X1 port map( A1 => n11792, A2 => n8432, B1 => n11788, B2 => 
                           n8656, ZN => n9856);
   U9845 : AOI221_X1 port map( B1 => n10975, B2 => n11800, C1 => n11167, C2 => 
                           n11796, A => n9839, ZN => n9836);
   U9846 : OAI22_X1 port map( A1 => n11792, A2 => n8431, B1 => n11788, B2 => 
                           n8655, ZN => n9839);
   U9847 : AOI221_X1 port map( B1 => n10976, B2 => n11800, C1 => n11168, C2 => 
                           n11796, A => n9822, ZN => n9819);
   U9848 : OAI22_X1 port map( A1 => n11792, A2 => n8430, B1 => n11788, B2 => 
                           n8654, ZN => n9822);
   U9849 : AOI221_X1 port map( B1 => n10977, B2 => n11800, C1 => n11169, C2 => 
                           n11796, A => n9805, ZN => n9802);
   U9850 : OAI22_X1 port map( A1 => n11792, A2 => n8429, B1 => n11788, B2 => 
                           n8653, ZN => n9805);
   U9851 : AOI221_X1 port map( B1 => n10978, B2 => n11800, C1 => n11170, C2 => 
                           n11796, A => n9788, ZN => n9785);
   U9852 : OAI22_X1 port map( A1 => n11792, A2 => n8428, B1 => n11788, B2 => 
                           n8652, ZN => n9788);
   U9853 : AOI221_X1 port map( B1 => n10979, B2 => n11800, C1 => n11171, C2 => 
                           n11796, A => n9771, ZN => n9768);
   U9854 : OAI22_X1 port map( A1 => n11792, A2 => n8427, B1 => n11788, B2 => 
                           n8651, ZN => n9771);
   U9855 : AOI221_X1 port map( B1 => n10980, B2 => n11800, C1 => n11172, C2 => 
                           n11796, A => n9754, ZN => n9751);
   U9856 : OAI22_X1 port map( A1 => n11792, A2 => n8426, B1 => n11788, B2 => 
                           n8650, ZN => n9754);
   U9857 : AOI221_X1 port map( B1 => n10981, B2 => n11800, C1 => n11173, C2 => 
                           n11796, A => n9737, ZN => n9734);
   U9858 : OAI22_X1 port map( A1 => n11792, A2 => n8425, B1 => n11788, B2 => 
                           n8649, ZN => n9737);
   U9859 : AOI221_X1 port map( B1 => n10982, B2 => n11800, C1 => n11174, C2 => 
                           n11796, A => n9720, ZN => n9717);
   U9860 : OAI22_X1 port map( A1 => n11792, A2 => n8424, B1 => n11788, B2 => 
                           n8648, ZN => n9720);
   U9861 : AOI221_X1 port map( B1 => n10983, B2 => n11800, C1 => n11175, C2 => 
                           n11796, A => n9703, ZN => n9700);
   U9862 : OAI22_X1 port map( A1 => n11792, A2 => n8423, B1 => n11788, B2 => 
                           n8647, ZN => n9703);
   U9863 : AOI221_X1 port map( B1 => n10984, B2 => n11800, C1 => n11176, C2 => 
                           n11796, A => n9686, ZN => n9683);
   U9864 : OAI22_X1 port map( A1 => n11792, A2 => n8422, B1 => n11788, B2 => 
                           n8646, ZN => n9686);
   U9865 : AOI221_X1 port map( B1 => n10985, B2 => n11801, C1 => n11177, C2 => 
                           n11797, A => n9669, ZN => n9666);
   U9866 : OAI22_X1 port map( A1 => n11793, A2 => n8421, B1 => n11789, B2 => 
                           n8645, ZN => n9669);
   U9867 : AOI221_X1 port map( B1 => n10986, B2 => n11801, C1 => n11178, C2 => 
                           n11797, A => n9652, ZN => n9649);
   U9868 : OAI22_X1 port map( A1 => n11793, A2 => n8420, B1 => n11789, B2 => 
                           n8644, ZN => n9652);
   U9869 : AOI221_X1 port map( B1 => n10987, B2 => n11801, C1 => n11179, C2 => 
                           n11797, A => n9635, ZN => n9632);
   U9870 : OAI22_X1 port map( A1 => n11793, A2 => n8419, B1 => n11789, B2 => 
                           n8643, ZN => n9635);
   U9871 : AOI221_X1 port map( B1 => n10988, B2 => n11801, C1 => n11180, C2 => 
                           n11797, A => n9618, ZN => n9615);
   U9872 : OAI22_X1 port map( A1 => n11793, A2 => n8418, B1 => n11789, B2 => 
                           n8642, ZN => n9618);
   U9873 : AOI221_X1 port map( B1 => n10989, B2 => n11801, C1 => n11181, C2 => 
                           n11797, A => n9601, ZN => n9598);
   U9874 : OAI22_X1 port map( A1 => n11793, A2 => n8417, B1 => n11789, B2 => 
                           n8641, ZN => n9601);
   U9875 : AOI221_X1 port map( B1 => n10990, B2 => n11801, C1 => n11182, C2 => 
                           n11797, A => n9584, ZN => n9581);
   U9876 : OAI22_X1 port map( A1 => n11793, A2 => n8416, B1 => n11789, B2 => 
                           n8640, ZN => n9584);
   U9877 : AOI221_X1 port map( B1 => n10991, B2 => n11801, C1 => n11183, C2 => 
                           n11797, A => n9567, ZN => n9564);
   U9878 : OAI22_X1 port map( A1 => n11793, A2 => n8415, B1 => n11789, B2 => 
                           n8639, ZN => n9567);
   U9879 : AOI221_X1 port map( B1 => n10992, B2 => n11801, C1 => n11184, C2 => 
                           n11797, A => n9550, ZN => n9547);
   U9880 : OAI22_X1 port map( A1 => n11793, A2 => n8414, B1 => n11789, B2 => 
                           n8638, ZN => n9550);
   U9881 : AOI221_X1 port map( B1 => n10993, B2 => n11801, C1 => n11185, C2 => 
                           n11797, A => n9533, ZN => n9530);
   U9882 : OAI22_X1 port map( A1 => n11793, A2 => n8413, B1 => n11789, B2 => 
                           n8637, ZN => n9533);
   U9883 : AOI221_X1 port map( B1 => n10994, B2 => n11801, C1 => n11186, C2 => 
                           n11797, A => n9516, ZN => n9513);
   U9884 : OAI22_X1 port map( A1 => n11793, A2 => n8412, B1 => n11789, B2 => 
                           n8636, ZN => n9516);
   U9885 : AOI221_X1 port map( B1 => n10995, B2 => n11801, C1 => n11187, C2 => 
                           n11797, A => n9499, ZN => n9496);
   U9886 : OAI22_X1 port map( A1 => n11793, A2 => n8411, B1 => n11789, B2 => 
                           n8635, ZN => n9499);
   U9887 : AOI221_X1 port map( B1 => n10996, B2 => n11801, C1 => n11188, C2 => 
                           n11797, A => n9482, ZN => n9479);
   U9888 : OAI22_X1 port map( A1 => n11793, A2 => n8410, B1 => n11789, B2 => 
                           n8634, ZN => n9482);
   U9889 : AOI221_X1 port map( B1 => n10997, B2 => n11802, C1 => n11189, C2 => 
                           n11798, A => n9465, ZN => n9462);
   U9890 : OAI22_X1 port map( A1 => n11794, A2 => n8409, B1 => n11790, B2 => 
                           n8633, ZN => n9465);
   U9891 : AOI221_X1 port map( B1 => n10998, B2 => n11802, C1 => n11190, C2 => 
                           n11798, A => n9448, ZN => n9445);
   U9892 : OAI22_X1 port map( A1 => n11794, A2 => n8408, B1 => n11790, B2 => 
                           n8632, ZN => n9448);
   U9893 : AOI221_X1 port map( B1 => n10999, B2 => n11802, C1 => n11191, C2 => 
                           n11798, A => n9431, ZN => n9428);
   U9894 : OAI22_X1 port map( A1 => n11794, A2 => n8407, B1 => n11790, B2 => 
                           n8631, ZN => n9431);
   U9895 : AOI221_X1 port map( B1 => n11000, B2 => n11802, C1 => n11192, C2 => 
                           n11798, A => n9414, ZN => n9411);
   U9896 : OAI22_X1 port map( A1 => n11794, A2 => n8406, B1 => n11790, B2 => 
                           n8630, ZN => n9414);
   U9897 : AOI221_X1 port map( B1 => n11001, B2 => n11802, C1 => n11193, C2 => 
                           n11798, A => n9397, ZN => n9394);
   U9898 : OAI22_X1 port map( A1 => n11794, A2 => n8405, B1 => n11790, B2 => 
                           n8629, ZN => n9397);
   U9899 : AOI221_X1 port map( B1 => n11002, B2 => n11802, C1 => n11194, C2 => 
                           n11798, A => n9380, ZN => n9377);
   U9900 : OAI22_X1 port map( A1 => n11794, A2 => n8404, B1 => n11790, B2 => 
                           n8628, ZN => n9380);
   U9901 : AOI221_X1 port map( B1 => n11003, B2 => n11802, C1 => n11195, C2 => 
                           n11798, A => n9363, ZN => n9360);
   U9902 : OAI22_X1 port map( A1 => n11794, A2 => n8403, B1 => n11790, B2 => 
                           n8627, ZN => n9363);
   U9903 : AOI221_X1 port map( B1 => n11004, B2 => n11802, C1 => n11196, C2 => 
                           n11798, A => n9335, ZN => n9325);
   U9904 : OAI22_X1 port map( A1 => n11794, A2 => n8402, B1 => n11790, B2 => 
                           n8626, ZN => n9335);
   U9905 : AOI221_X1 port map( B1 => n11663, B2 => n10997, C1 => n11659, C2 => 
                           n11189, A => n10055, ZN => n10052);
   U9906 : OAI22_X1 port map( A1 => n8409, A2 => n11655, B1 => n8633, B2 => 
                           n11651, ZN => n10055);
   U9907 : AOI221_X1 port map( B1 => n11663, B2 => n10998, C1 => n11659, C2 => 
                           n11190, A => n10038, ZN => n10035);
   U9908 : OAI22_X1 port map( A1 => n8408, A2 => n11655, B1 => n8632, B2 => 
                           n11651, ZN => n10038);
   U9909 : AOI221_X1 port map( B1 => n11663, B2 => n10999, C1 => n11659, C2 => 
                           n11191, A => n10021, ZN => n10018);
   U9910 : OAI22_X1 port map( A1 => n8407, A2 => n11655, B1 => n8631, B2 => 
                           n11651, ZN => n10021);
   U9911 : AOI221_X1 port map( B1 => n11663, B2 => n11000, C1 => n11659, C2 => 
                           n11192, A => n10004, ZN => n10001);
   U9912 : OAI22_X1 port map( A1 => n8406, A2 => n11655, B1 => n8630, B2 => 
                           n11651, ZN => n10004);
   U9913 : AOI221_X1 port map( B1 => n11663, B2 => n11001, C1 => n11659, C2 => 
                           n11193, A => n9987, ZN => n9984);
   U9914 : OAI22_X1 port map( A1 => n8405, A2 => n11655, B1 => n8629, B2 => 
                           n11651, ZN => n9987);
   U9915 : AOI221_X1 port map( B1 => n11663, B2 => n11002, C1 => n11659, C2 => 
                           n11194, A => n9970, ZN => n9967);
   U9916 : OAI22_X1 port map( A1 => n8404, A2 => n11655, B1 => n8628, B2 => 
                           n11651, ZN => n9970);
   U9917 : AOI221_X1 port map( B1 => n11663, B2 => n11003, C1 => n11659, C2 => 
                           n11195, A => n9953, ZN => n9950);
   U9918 : OAI22_X1 port map( A1 => n8403, A2 => n11655, B1 => n8627, B2 => 
                           n11651, ZN => n9953);
   U9919 : AOI221_X1 port map( B1 => n11663, B2 => n11004, C1 => n11659, C2 => 
                           n11196, A => n9925, ZN => n9915);
   U9920 : OAI22_X1 port map( A1 => n8402, A2 => n11655, B1 => n8626, B2 => 
                           n11651, ZN => n9925);
   U9921 : AOI221_X1 port map( B1 => n11661, B2 => n10973, C1 => n11657, C2 => 
                           n11165, A => n10475, ZN => n10469);
   U9922 : OAI22_X1 port map( A1 => n8433, A2 => n11653, B1 => n8657, B2 => 
                           n11649, ZN => n10475);
   U9923 : AOI221_X1 port map( B1 => n11661, B2 => n10974, C1 => n11657, C2 => 
                           n11166, A => n10446, ZN => n10443);
   U9924 : OAI22_X1 port map( A1 => n8432, A2 => n11653, B1 => n8656, B2 => 
                           n11649, ZN => n10446);
   U9925 : AOI221_X1 port map( B1 => n11661, B2 => n10975, C1 => n11657, C2 => 
                           n11167, A => n10429, ZN => n10426);
   U9926 : OAI22_X1 port map( A1 => n8431, A2 => n11653, B1 => n8655, B2 => 
                           n11649, ZN => n10429);
   U9927 : AOI221_X1 port map( B1 => n11661, B2 => n10976, C1 => n11657, C2 => 
                           n11168, A => n10412, ZN => n10409);
   U9928 : OAI22_X1 port map( A1 => n8430, A2 => n11653, B1 => n8654, B2 => 
                           n11649, ZN => n10412);
   U9929 : AOI221_X1 port map( B1 => n11661, B2 => n10977, C1 => n11657, C2 => 
                           n11169, A => n10395, ZN => n10392);
   U9930 : OAI22_X1 port map( A1 => n8429, A2 => n11653, B1 => n8653, B2 => 
                           n11649, ZN => n10395);
   U9931 : AOI221_X1 port map( B1 => n11661, B2 => n10978, C1 => n11657, C2 => 
                           n11170, A => n10378, ZN => n10375);
   U9932 : OAI22_X1 port map( A1 => n8428, A2 => n11653, B1 => n8652, B2 => 
                           n11649, ZN => n10378);
   U9933 : AOI221_X1 port map( B1 => n11661, B2 => n10979, C1 => n11657, C2 => 
                           n11171, A => n10361, ZN => n10358);
   U9934 : OAI22_X1 port map( A1 => n8427, A2 => n11653, B1 => n8651, B2 => 
                           n11649, ZN => n10361);
   U9935 : AOI221_X1 port map( B1 => n11661, B2 => n10980, C1 => n11657, C2 => 
                           n11172, A => n10344, ZN => n10341);
   U9936 : OAI22_X1 port map( A1 => n8426, A2 => n11653, B1 => n8650, B2 => 
                           n11649, ZN => n10344);
   U9937 : AOI221_X1 port map( B1 => n11661, B2 => n10981, C1 => n11657, C2 => 
                           n11173, A => n10327, ZN => n10324);
   U9938 : OAI22_X1 port map( A1 => n8425, A2 => n11653, B1 => n8649, B2 => 
                           n11649, ZN => n10327);
   U9939 : AOI221_X1 port map( B1 => n11661, B2 => n10982, C1 => n11657, C2 => 
                           n11174, A => n10310, ZN => n10307);
   U9940 : OAI22_X1 port map( A1 => n8424, A2 => n11653, B1 => n8648, B2 => 
                           n11649, ZN => n10310);
   U9941 : AOI221_X1 port map( B1 => n11661, B2 => n10983, C1 => n11657, C2 => 
                           n11175, A => n10293, ZN => n10290);
   U9942 : OAI22_X1 port map( A1 => n8423, A2 => n11653, B1 => n8647, B2 => 
                           n11649, ZN => n10293);
   U9943 : AOI221_X1 port map( B1 => n11661, B2 => n10984, C1 => n11657, C2 => 
                           n11176, A => n10276, ZN => n10273);
   U9944 : OAI22_X1 port map( A1 => n8422, A2 => n11653, B1 => n8646, B2 => 
                           n11649, ZN => n10276);
   U9945 : AOI221_X1 port map( B1 => n11662, B2 => n10985, C1 => n11658, C2 => 
                           n11177, A => n10259, ZN => n10256);
   U9946 : OAI22_X1 port map( A1 => n8421, A2 => n11654, B1 => n8645, B2 => 
                           n11650, ZN => n10259);
   U9947 : AOI221_X1 port map( B1 => n11662, B2 => n10986, C1 => n11658, C2 => 
                           n11178, A => n10242, ZN => n10239);
   U9948 : OAI22_X1 port map( A1 => n8420, A2 => n11654, B1 => n8644, B2 => 
                           n11650, ZN => n10242);
   U9949 : AOI221_X1 port map( B1 => n11662, B2 => n10987, C1 => n11658, C2 => 
                           n11179, A => n10225, ZN => n10222);
   U9950 : OAI22_X1 port map( A1 => n8419, A2 => n11654, B1 => n8643, B2 => 
                           n11650, ZN => n10225);
   U9951 : AOI221_X1 port map( B1 => n11662, B2 => n10988, C1 => n11658, C2 => 
                           n11180, A => n10208, ZN => n10205);
   U9952 : OAI22_X1 port map( A1 => n8418, A2 => n11654, B1 => n8642, B2 => 
                           n11650, ZN => n10208);
   U9953 : AOI221_X1 port map( B1 => n11662, B2 => n10989, C1 => n11658, C2 => 
                           n11181, A => n10191, ZN => n10188);
   U9954 : OAI22_X1 port map( A1 => n8417, A2 => n11654, B1 => n8641, B2 => 
                           n11650, ZN => n10191);
   U9955 : AOI221_X1 port map( B1 => n11662, B2 => n10990, C1 => n11658, C2 => 
                           n11182, A => n10174, ZN => n10171);
   U9956 : OAI22_X1 port map( A1 => n8416, A2 => n11654, B1 => n8640, B2 => 
                           n11650, ZN => n10174);
   U9957 : AOI221_X1 port map( B1 => n11662, B2 => n10991, C1 => n11658, C2 => 
                           n11183, A => n10157, ZN => n10154);
   U9958 : OAI22_X1 port map( A1 => n8415, A2 => n11654, B1 => n8639, B2 => 
                           n11650, ZN => n10157);
   U9959 : AOI221_X1 port map( B1 => n11662, B2 => n10992, C1 => n11658, C2 => 
                           n11184, A => n10140, ZN => n10137);
   U9960 : OAI22_X1 port map( A1 => n8414, A2 => n11654, B1 => n8638, B2 => 
                           n11650, ZN => n10140);
   U9961 : AOI221_X1 port map( B1 => n11662, B2 => n10993, C1 => n11658, C2 => 
                           n11185, A => n10123, ZN => n10120);
   U9962 : OAI22_X1 port map( A1 => n8413, A2 => n11654, B1 => n8637, B2 => 
                           n11650, ZN => n10123);
   U9963 : AOI221_X1 port map( B1 => n11662, B2 => n10994, C1 => n11658, C2 => 
                           n11186, A => n10106, ZN => n10103);
   U9964 : OAI22_X1 port map( A1 => n8412, A2 => n11654, B1 => n8636, B2 => 
                           n11650, ZN => n10106);
   U9965 : AOI221_X1 port map( B1 => n11662, B2 => n10995, C1 => n11658, C2 => 
                           n11187, A => n10089, ZN => n10086);
   U9966 : OAI22_X1 port map( A1 => n8411, A2 => n11654, B1 => n8635, B2 => 
                           n11650, ZN => n10089);
   U9967 : AOI221_X1 port map( B1 => n11662, B2 => n10996, C1 => n11658, C2 => 
                           n11188, A => n10072, ZN => n10069);
   U9968 : OAI22_X1 port map( A1 => n8410, A2 => n11654, B1 => n8634, B2 => 
                           n11650, ZN => n10072);
   U9969 : OAI22_X1 port map( A1 => n11274, A2 => n11483, B1 => n9169, B2 => 
                           n11372, ZN => n1406);
   U9970 : OAI22_X1 port map( A1 => n11274, A2 => n11487, B1 => n9168, B2 => 
                           n11372, ZN => n1407);
   U9971 : OAI22_X1 port map( A1 => n11274, A2 => n11491, B1 => n9167, B2 => 
                           n11372, ZN => n1408);
   U9972 : OAI22_X1 port map( A1 => n11274, A2 => n11495, B1 => n9166, B2 => 
                           n11372, ZN => n1409);
   U9973 : OAI22_X1 port map( A1 => n11274, A2 => n11499, B1 => n9165, B2 => 
                           n11372, ZN => n1410);
   U9974 : OAI22_X1 port map( A1 => n11274, A2 => n11503, B1 => n9164, B2 => 
                           n11372, ZN => n1411);
   U9975 : OAI22_X1 port map( A1 => n11274, A2 => n11507, B1 => n9163, B2 => 
                           n11372, ZN => n1412);
   U9976 : OAI22_X1 port map( A1 => n11274, A2 => n11511, B1 => n9162, B2 => 
                           n11372, ZN => n1413);
   U9977 : OAI22_X1 port map( A1 => n11273, A2 => n11515, B1 => n9161, B2 => 
                           n11372, ZN => n1414);
   U9978 : OAI22_X1 port map( A1 => n11273, A2 => n11519, B1 => n9160, B2 => 
                           n11372, ZN => n1415);
   U9979 : OAI22_X1 port map( A1 => n11273, A2 => n11523, B1 => n9159, B2 => 
                           n11372, ZN => n1416);
   U9980 : OAI22_X1 port map( A1 => n11273, A2 => n11527, B1 => n9158, B2 => 
                           n11372, ZN => n1417);
   U9981 : OAI22_X1 port map( A1 => n11273, A2 => n11531, B1 => n9157, B2 => 
                           n10550, ZN => n1418);
   U9982 : OAI22_X1 port map( A1 => n11273, A2 => n11535, B1 => n9156, B2 => 
                           n10550, ZN => n1419);
   U9983 : OAI22_X1 port map( A1 => n11273, A2 => n11539, B1 => n9155, B2 => 
                           n10550, ZN => n1420);
   U9984 : OAI22_X1 port map( A1 => n11273, A2 => n11543, B1 => n9154, B2 => 
                           n11372, ZN => n1421);
   U9985 : OAI22_X1 port map( A1 => n11273, A2 => n11547, B1 => n9153, B2 => 
                           n11372, ZN => n1422);
   U9986 : OAI22_X1 port map( A1 => n11273, A2 => n11551, B1 => n9152, B2 => 
                           n11372, ZN => n1423);
   U9987 : OAI22_X1 port map( A1 => n11273, A2 => n11555, B1 => n9151, B2 => 
                           n11372, ZN => n1424);
   U9988 : OAI22_X1 port map( A1 => n11273, A2 => n11559, B1 => n9150, B2 => 
                           n11372, ZN => n1425);
   U9989 : OAI22_X1 port map( A1 => n11272, A2 => n11563, B1 => n9149, B2 => 
                           n11372, ZN => n1426);
   U9990 : OAI22_X1 port map( A1 => n11272, A2 => n11567, B1 => n9148, B2 => 
                           n11372, ZN => n1427);
   U9991 : OAI22_X1 port map( A1 => n11272, A2 => n11571, B1 => n9147, B2 => 
                           n11372, ZN => n1428);
   U9992 : OAI22_X1 port map( A1 => n11272, A2 => n11575, B1 => n9146, B2 => 
                           n11372, ZN => n1429);
   U9993 : OAI22_X1 port map( A1 => n11272, A2 => n11579, B1 => n9145, B2 => 
                           n10550, ZN => n1430);
   U9994 : OAI22_X1 port map( A1 => n11272, A2 => n11583, B1 => n9144, B2 => 
                           n10550, ZN => n1431);
   U9995 : OAI22_X1 port map( A1 => n11272, A2 => n11587, B1 => n9143, B2 => 
                           n10550, ZN => n1432);
   U9996 : OAI22_X1 port map( A1 => n11272, A2 => n11591, B1 => n9142, B2 => 
                           n10550, ZN => n1433);
   U9997 : OAI22_X1 port map( A1 => n11272, A2 => n11595, B1 => n9141, B2 => 
                           n10550, ZN => n1434);
   U9998 : OAI22_X1 port map( A1 => n11272, A2 => n11599, B1 => n9140, B2 => 
                           n10550, ZN => n1435);
   U9999 : OAI22_X1 port map( A1 => n11272, A2 => n11603, B1 => n9139, B2 => 
                           n10550, ZN => n1436);
   U10000 : OAI22_X1 port map( A1 => n11272, A2 => n11611, B1 => n9138, B2 => 
                           n10550, ZN => n1437);
   U10001 : OAI22_X1 port map( A1 => n11283, A2 => n11483, B1 => n9073, B2 => 
                           n11384, ZN => n1502);
   U10002 : OAI22_X1 port map( A1 => n11283, A2 => n11487, B1 => n9072, B2 => 
                           n11384, ZN => n1503);
   U10003 : OAI22_X1 port map( A1 => n11283, A2 => n11491, B1 => n9071, B2 => 
                           n11384, ZN => n1504);
   U10004 : OAI22_X1 port map( A1 => n11283, A2 => n11495, B1 => n9070, B2 => 
                           n11384, ZN => n1505);
   U10005 : OAI22_X1 port map( A1 => n11283, A2 => n11499, B1 => n9069, B2 => 
                           n11384, ZN => n1506);
   U10006 : OAI22_X1 port map( A1 => n11283, A2 => n11503, B1 => n9068, B2 => 
                           n11384, ZN => n1507);
   U10007 : OAI22_X1 port map( A1 => n11283, A2 => n11507, B1 => n9067, B2 => 
                           n11384, ZN => n1508);
   U10008 : OAI22_X1 port map( A1 => n11283, A2 => n11511, B1 => n9066, B2 => 
                           n11384, ZN => n1509);
   U10009 : OAI22_X1 port map( A1 => n11282, A2 => n11515, B1 => n9065, B2 => 
                           n11384, ZN => n1510);
   U10010 : OAI22_X1 port map( A1 => n11282, A2 => n11519, B1 => n9064, B2 => 
                           n11384, ZN => n1511);
   U10011 : OAI22_X1 port map( A1 => n11282, A2 => n11523, B1 => n9063, B2 => 
                           n11384, ZN => n1512);
   U10012 : OAI22_X1 port map( A1 => n11282, A2 => n11527, B1 => n9062, B2 => 
                           n11384, ZN => n1513);
   U10013 : OAI22_X1 port map( A1 => n11282, A2 => n11531, B1 => n9061, B2 => 
                           n10546, ZN => n1514);
   U10014 : OAI22_X1 port map( A1 => n11282, A2 => n11535, B1 => n9060, B2 => 
                           n10546, ZN => n1515);
   U10015 : OAI22_X1 port map( A1 => n11282, A2 => n11539, B1 => n9059, B2 => 
                           n10546, ZN => n1516);
   U10016 : OAI22_X1 port map( A1 => n11282, A2 => n11543, B1 => n9058, B2 => 
                           n11384, ZN => n1517);
   U10017 : OAI22_X1 port map( A1 => n11282, A2 => n11547, B1 => n9057, B2 => 
                           n11384, ZN => n1518);
   U10018 : OAI22_X1 port map( A1 => n11282, A2 => n11551, B1 => n9056, B2 => 
                           n11384, ZN => n1519);
   U10019 : OAI22_X1 port map( A1 => n11282, A2 => n11555, B1 => n9055, B2 => 
                           n11384, ZN => n1520);
   U10020 : OAI22_X1 port map( A1 => n11282, A2 => n11559, B1 => n9054, B2 => 
                           n11384, ZN => n1521);
   U10021 : OAI22_X1 port map( A1 => n11281, A2 => n11563, B1 => n9053, B2 => 
                           n11384, ZN => n1522);
   U10022 : OAI22_X1 port map( A1 => n11281, A2 => n11567, B1 => n9052, B2 => 
                           n11384, ZN => n1523);
   U10023 : OAI22_X1 port map( A1 => n11281, A2 => n11571, B1 => n9051, B2 => 
                           n11384, ZN => n1524);
   U10024 : OAI22_X1 port map( A1 => n11281, A2 => n11575, B1 => n9050, B2 => 
                           n11384, ZN => n1525);
   U10025 : OAI22_X1 port map( A1 => n11281, A2 => n11579, B1 => n9049, B2 => 
                           n10546, ZN => n1526);
   U10026 : OAI22_X1 port map( A1 => n11281, A2 => n11583, B1 => n9048, B2 => 
                           n10546, ZN => n1527);
   U10027 : OAI22_X1 port map( A1 => n11281, A2 => n11587, B1 => n9047, B2 => 
                           n10546, ZN => n1528);
   U10028 : OAI22_X1 port map( A1 => n11281, A2 => n11591, B1 => n9046, B2 => 
                           n10546, ZN => n1529);
   U10029 : OAI22_X1 port map( A1 => n11281, A2 => n11595, B1 => n9045, B2 => 
                           n10546, ZN => n1530);
   U10030 : OAI22_X1 port map( A1 => n11281, A2 => n11599, B1 => n9044, B2 => 
                           n10546, ZN => n1531);
   U10031 : OAI22_X1 port map( A1 => n11281, A2 => n11603, B1 => n9043, B2 => 
                           n10546, ZN => n1532);
   U10032 : OAI22_X1 port map( A1 => n11281, A2 => n11611, B1 => n9042, B2 => 
                           n10546, ZN => n1533);
   U10033 : OAI22_X1 port map( A1 => n11286, A2 => n11482, B1 => n9041, B2 => 
                           n11388, ZN => n1534);
   U10034 : OAI22_X1 port map( A1 => n11286, A2 => n11486, B1 => n9040, B2 => 
                           n11388, ZN => n1535);
   U10035 : OAI22_X1 port map( A1 => n11286, A2 => n11490, B1 => n9039, B2 => 
                           n11388, ZN => n1536);
   U10036 : OAI22_X1 port map( A1 => n11286, A2 => n11494, B1 => n9038, B2 => 
                           n11388, ZN => n1537);
   U10037 : OAI22_X1 port map( A1 => n11286, A2 => n11498, B1 => n9037, B2 => 
                           n11388, ZN => n1538);
   U10038 : OAI22_X1 port map( A1 => n11286, A2 => n11502, B1 => n9036, B2 => 
                           n11388, ZN => n1539);
   U10039 : OAI22_X1 port map( A1 => n11286, A2 => n11506, B1 => n9035, B2 => 
                           n11388, ZN => n1540);
   U10040 : OAI22_X1 port map( A1 => n11286, A2 => n11510, B1 => n9034, B2 => 
                           n11388, ZN => n1541);
   U10041 : OAI22_X1 port map( A1 => n11285, A2 => n11514, B1 => n9033, B2 => 
                           n11388, ZN => n1542);
   U10042 : OAI22_X1 port map( A1 => n11285, A2 => n11518, B1 => n9032, B2 => 
                           n11388, ZN => n1543);
   U10043 : OAI22_X1 port map( A1 => n11285, A2 => n11522, B1 => n9031, B2 => 
                           n11388, ZN => n1544);
   U10044 : OAI22_X1 port map( A1 => n11285, A2 => n11526, B1 => n9030, B2 => 
                           n11388, ZN => n1545);
   U10045 : OAI22_X1 port map( A1 => n11285, A2 => n11530, B1 => n9029, B2 => 
                           n10545, ZN => n1546);
   U10046 : OAI22_X1 port map( A1 => n11285, A2 => n11534, B1 => n9028, B2 => 
                           n10545, ZN => n1547);
   U10047 : OAI22_X1 port map( A1 => n11285, A2 => n11538, B1 => n9027, B2 => 
                           n10545, ZN => n1548);
   U10048 : OAI22_X1 port map( A1 => n11285, A2 => n11542, B1 => n9026, B2 => 
                           n11388, ZN => n1549);
   U10049 : OAI22_X1 port map( A1 => n11285, A2 => n11546, B1 => n9025, B2 => 
                           n11388, ZN => n1550);
   U10050 : OAI22_X1 port map( A1 => n11285, A2 => n11550, B1 => n9024, B2 => 
                           n11388, ZN => n1551);
   U10051 : OAI22_X1 port map( A1 => n11285, A2 => n11554, B1 => n9023, B2 => 
                           n11388, ZN => n1552);
   U10052 : OAI22_X1 port map( A1 => n11285, A2 => n11558, B1 => n9022, B2 => 
                           n11388, ZN => n1553);
   U10053 : OAI22_X1 port map( A1 => n11284, A2 => n11562, B1 => n9021, B2 => 
                           n11388, ZN => n1554);
   U10054 : OAI22_X1 port map( A1 => n11284, A2 => n11566, B1 => n9020, B2 => 
                           n11388, ZN => n1555);
   U10055 : OAI22_X1 port map( A1 => n11284, A2 => n11570, B1 => n9019, B2 => 
                           n11388, ZN => n1556);
   U10056 : OAI22_X1 port map( A1 => n11284, A2 => n11574, B1 => n9018, B2 => 
                           n11388, ZN => n1557);
   U10057 : OAI22_X1 port map( A1 => n11284, A2 => n11578, B1 => n9017, B2 => 
                           n10545, ZN => n1558);
   U10058 : OAI22_X1 port map( A1 => n11284, A2 => n11582, B1 => n9016, B2 => 
                           n10545, ZN => n1559);
   U10059 : OAI22_X1 port map( A1 => n11284, A2 => n11586, B1 => n9015, B2 => 
                           n10545, ZN => n1560);
   U10060 : OAI22_X1 port map( A1 => n11284, A2 => n11590, B1 => n9014, B2 => 
                           n10545, ZN => n1561);
   U10061 : OAI22_X1 port map( A1 => n11284, A2 => n11594, B1 => n9013, B2 => 
                           n10545, ZN => n1562);
   U10062 : OAI22_X1 port map( A1 => n11284, A2 => n11598, B1 => n9012, B2 => 
                           n10545, ZN => n1563);
   U10063 : OAI22_X1 port map( A1 => n11284, A2 => n11602, B1 => n9011, B2 => 
                           n10545, ZN => n1564);
   U10064 : OAI22_X1 port map( A1 => n11284, A2 => n11610, B1 => n9010, B2 => 
                           n10545, ZN => n1565);
   U10065 : OAI22_X1 port map( A1 => n11313, A2 => n11482, B1 => n8753, B2 => 
                           n11424, ZN => n1822);
   U10066 : OAI22_X1 port map( A1 => n11313, A2 => n11486, B1 => n8752, B2 => 
                           n11424, ZN => n1823);
   U10067 : OAI22_X1 port map( A1 => n11313, A2 => n11490, B1 => n8751, B2 => 
                           n11424, ZN => n1824);
   U10068 : OAI22_X1 port map( A1 => n11313, A2 => n11494, B1 => n8750, B2 => 
                           n11424, ZN => n1825);
   U10069 : OAI22_X1 port map( A1 => n11313, A2 => n11498, B1 => n8749, B2 => 
                           n11424, ZN => n1826);
   U10070 : OAI22_X1 port map( A1 => n11313, A2 => n11502, B1 => n8748, B2 => 
                           n11424, ZN => n1827);
   U10071 : OAI22_X1 port map( A1 => n11313, A2 => n11506, B1 => n8747, B2 => 
                           n11424, ZN => n1828);
   U10072 : OAI22_X1 port map( A1 => n11313, A2 => n11510, B1 => n8746, B2 => 
                           n11424, ZN => n1829);
   U10073 : OAI22_X1 port map( A1 => n11312, A2 => n11514, B1 => n8745, B2 => 
                           n11424, ZN => n1830);
   U10074 : OAI22_X1 port map( A1 => n11312, A2 => n11518, B1 => n8744, B2 => 
                           n11424, ZN => n1831);
   U10075 : OAI22_X1 port map( A1 => n11312, A2 => n11522, B1 => n8743, B2 => 
                           n11424, ZN => n1832);
   U10076 : OAI22_X1 port map( A1 => n11312, A2 => n11526, B1 => n8742, B2 => 
                           n11424, ZN => n1833);
   U10077 : OAI22_X1 port map( A1 => n11312, A2 => n11530, B1 => n8741, B2 => 
                           n10533, ZN => n1834);
   U10078 : OAI22_X1 port map( A1 => n11312, A2 => n11534, B1 => n8740, B2 => 
                           n10533, ZN => n1835);
   U10079 : OAI22_X1 port map( A1 => n11312, A2 => n11538, B1 => n8739, B2 => 
                           n10533, ZN => n1836);
   U10080 : OAI22_X1 port map( A1 => n11312, A2 => n11542, B1 => n8738, B2 => 
                           n11424, ZN => n1837);
   U10081 : OAI22_X1 port map( A1 => n11312, A2 => n11546, B1 => n8737, B2 => 
                           n11424, ZN => n1838);
   U10082 : OAI22_X1 port map( A1 => n11312, A2 => n11550, B1 => n8736, B2 => 
                           n11424, ZN => n1839);
   U10083 : OAI22_X1 port map( A1 => n11312, A2 => n11554, B1 => n8735, B2 => 
                           n11424, ZN => n1840);
   U10084 : OAI22_X1 port map( A1 => n11312, A2 => n11558, B1 => n8734, B2 => 
                           n11424, ZN => n1841);
   U10085 : OAI22_X1 port map( A1 => n11311, A2 => n11562, B1 => n8733, B2 => 
                           n11424, ZN => n1842);
   U10086 : OAI22_X1 port map( A1 => n11311, A2 => n11566, B1 => n8732, B2 => 
                           n11424, ZN => n1843);
   U10087 : OAI22_X1 port map( A1 => n11311, A2 => n11570, B1 => n8731, B2 => 
                           n11424, ZN => n1844);
   U10088 : OAI22_X1 port map( A1 => n11311, A2 => n11574, B1 => n8730, B2 => 
                           n11424, ZN => n1845);
   U10089 : OAI22_X1 port map( A1 => n11311, A2 => n11578, B1 => n8729, B2 => 
                           n10533, ZN => n1846);
   U10090 : OAI22_X1 port map( A1 => n11311, A2 => n11582, B1 => n8728, B2 => 
                           n10533, ZN => n1847);
   U10091 : OAI22_X1 port map( A1 => n11311, A2 => n11586, B1 => n8727, B2 => 
                           n10533, ZN => n1848);
   U10092 : OAI22_X1 port map( A1 => n11311, A2 => n11590, B1 => n8726, B2 => 
                           n10533, ZN => n1849);
   U10093 : OAI22_X1 port map( A1 => n11311, A2 => n11594, B1 => n8725, B2 => 
                           n10533, ZN => n1850);
   U10094 : OAI22_X1 port map( A1 => n11311, A2 => n11598, B1 => n8724, B2 => 
                           n10533, ZN => n1851);
   U10095 : OAI22_X1 port map( A1 => n11311, A2 => n11602, B1 => n8723, B2 => 
                           n10533, ZN => n1852);
   U10096 : OAI22_X1 port map( A1 => n11311, A2 => n11610, B1 => n8722, B2 => 
                           n10533, ZN => n1853);
   U10097 : OAI22_X1 port map( A1 => n11331, A2 => n11481, B1 => n8561, B2 => 
                           n11448, ZN => n2014);
   U10098 : OAI22_X1 port map( A1 => n11331, A2 => n11485, B1 => n8560, B2 => 
                           n11448, ZN => n2015);
   U10099 : OAI22_X1 port map( A1 => n11331, A2 => n11489, B1 => n8559, B2 => 
                           n11448, ZN => n2016);
   U10100 : OAI22_X1 port map( A1 => n11331, A2 => n11493, B1 => n8558, B2 => 
                           n11448, ZN => n2017);
   U10101 : OAI22_X1 port map( A1 => n11331, A2 => n11497, B1 => n8557, B2 => 
                           n11448, ZN => n2018);
   U10102 : OAI22_X1 port map( A1 => n11331, A2 => n11501, B1 => n8556, B2 => 
                           n11448, ZN => n2019);
   U10103 : OAI22_X1 port map( A1 => n11331, A2 => n11505, B1 => n8555, B2 => 
                           n11448, ZN => n2020);
   U10104 : OAI22_X1 port map( A1 => n11331, A2 => n11509, B1 => n8554, B2 => 
                           n11448, ZN => n2021);
   U10105 : OAI22_X1 port map( A1 => n11330, A2 => n11513, B1 => n8553, B2 => 
                           n11448, ZN => n2022);
   U10106 : OAI22_X1 port map( A1 => n11330, A2 => n11517, B1 => n8552, B2 => 
                           n11448, ZN => n2023);
   U10107 : OAI22_X1 port map( A1 => n11330, A2 => n11521, B1 => n8551, B2 => 
                           n11448, ZN => n2024);
   U10108 : OAI22_X1 port map( A1 => n11330, A2 => n11525, B1 => n8550, B2 => 
                           n11448, ZN => n2025);
   U10109 : OAI22_X1 port map( A1 => n11330, A2 => n11529, B1 => n8549, B2 => 
                           n10525, ZN => n2026);
   U10110 : OAI22_X1 port map( A1 => n11330, A2 => n11533, B1 => n8548, B2 => 
                           n10525, ZN => n2027);
   U10111 : OAI22_X1 port map( A1 => n11330, A2 => n11537, B1 => n8547, B2 => 
                           n10525, ZN => n2028);
   U10112 : OAI22_X1 port map( A1 => n11330, A2 => n11541, B1 => n8546, B2 => 
                           n11448, ZN => n2029);
   U10113 : OAI22_X1 port map( A1 => n11330, A2 => n11545, B1 => n8545, B2 => 
                           n11448, ZN => n2030);
   U10114 : OAI22_X1 port map( A1 => n11330, A2 => n11549, B1 => n8544, B2 => 
                           n11448, ZN => n2031);
   U10115 : OAI22_X1 port map( A1 => n11330, A2 => n11553, B1 => n8543, B2 => 
                           n11448, ZN => n2032);
   U10116 : OAI22_X1 port map( A1 => n11330, A2 => n11557, B1 => n8542, B2 => 
                           n11448, ZN => n2033);
   U10117 : OAI22_X1 port map( A1 => n11329, A2 => n11561, B1 => n8541, B2 => 
                           n11448, ZN => n2034);
   U10118 : OAI22_X1 port map( A1 => n11329, A2 => n11565, B1 => n8540, B2 => 
                           n11448, ZN => n2035);
   U10119 : OAI22_X1 port map( A1 => n11329, A2 => n11569, B1 => n8539, B2 => 
                           n11448, ZN => n2036);
   U10120 : OAI22_X1 port map( A1 => n11329, A2 => n11573, B1 => n8538, B2 => 
                           n11448, ZN => n2037);
   U10121 : OAI22_X1 port map( A1 => n11329, A2 => n11577, B1 => n8537, B2 => 
                           n10525, ZN => n2038);
   U10122 : OAI22_X1 port map( A1 => n11329, A2 => n11581, B1 => n8536, B2 => 
                           n10525, ZN => n2039);
   U10123 : OAI22_X1 port map( A1 => n11329, A2 => n11585, B1 => n8535, B2 => 
                           n10525, ZN => n2040);
   U10124 : OAI22_X1 port map( A1 => n11329, A2 => n11589, B1 => n8534, B2 => 
                           n10525, ZN => n2041);
   U10125 : OAI22_X1 port map( A1 => n11329, A2 => n11593, B1 => n8533, B2 => 
                           n10525, ZN => n2042);
   U10126 : OAI22_X1 port map( A1 => n11329, A2 => n11597, B1 => n8532, B2 => 
                           n10525, ZN => n2043);
   U10127 : OAI22_X1 port map( A1 => n11329, A2 => n11601, B1 => n8531, B2 => 
                           n10525, ZN => n2044);
   U10128 : OAI22_X1 port map( A1 => n11329, A2 => n11609, B1 => n8530, B2 => 
                           n10525, ZN => n2045);
   U10129 : OAI22_X1 port map( A1 => n11334, A2 => n11481, B1 => n8529, B2 => 
                           n11452, ZN => n2046);
   U10130 : OAI22_X1 port map( A1 => n11334, A2 => n11485, B1 => n8528, B2 => 
                           n11452, ZN => n2047);
   U10131 : OAI22_X1 port map( A1 => n11334, A2 => n11489, B1 => n8527, B2 => 
                           n11452, ZN => n2048);
   U10132 : OAI22_X1 port map( A1 => n11334, A2 => n11493, B1 => n8526, B2 => 
                           n11452, ZN => n2049);
   U10133 : OAI22_X1 port map( A1 => n11334, A2 => n11497, B1 => n8525, B2 => 
                           n11452, ZN => n2050);
   U10134 : OAI22_X1 port map( A1 => n11334, A2 => n11501, B1 => n8524, B2 => 
                           n11452, ZN => n2051);
   U10135 : OAI22_X1 port map( A1 => n11334, A2 => n11505, B1 => n8523, B2 => 
                           n11452, ZN => n2052);
   U10136 : OAI22_X1 port map( A1 => n11334, A2 => n11509, B1 => n8522, B2 => 
                           n11452, ZN => n2053);
   U10137 : OAI22_X1 port map( A1 => n11333, A2 => n11513, B1 => n8521, B2 => 
                           n11452, ZN => n2054);
   U10138 : OAI22_X1 port map( A1 => n11333, A2 => n11517, B1 => n8520, B2 => 
                           n11452, ZN => n2055);
   U10139 : OAI22_X1 port map( A1 => n11333, A2 => n11521, B1 => n8519, B2 => 
                           n11452, ZN => n2056);
   U10140 : OAI22_X1 port map( A1 => n11333, A2 => n11525, B1 => n8518, B2 => 
                           n11452, ZN => n2057);
   U10141 : OAI22_X1 port map( A1 => n11333, A2 => n11529, B1 => n8517, B2 => 
                           n10524, ZN => n2058);
   U10142 : OAI22_X1 port map( A1 => n11333, A2 => n11533, B1 => n8516, B2 => 
                           n10524, ZN => n2059);
   U10143 : OAI22_X1 port map( A1 => n11333, A2 => n11537, B1 => n8515, B2 => 
                           n10524, ZN => n2060);
   U10144 : OAI22_X1 port map( A1 => n11333, A2 => n11541, B1 => n8514, B2 => 
                           n11452, ZN => n2061);
   U10145 : OAI22_X1 port map( A1 => n11333, A2 => n11545, B1 => n8513, B2 => 
                           n11452, ZN => n2062);
   U10146 : OAI22_X1 port map( A1 => n11333, A2 => n11549, B1 => n8512, B2 => 
                           n11452, ZN => n2063);
   U10147 : OAI22_X1 port map( A1 => n11333, A2 => n11553, B1 => n8511, B2 => 
                           n11452, ZN => n2064);
   U10148 : OAI22_X1 port map( A1 => n11333, A2 => n11557, B1 => n8510, B2 => 
                           n11452, ZN => n2065);
   U10149 : OAI22_X1 port map( A1 => n11332, A2 => n11561, B1 => n8509, B2 => 
                           n11452, ZN => n2066);
   U10150 : OAI22_X1 port map( A1 => n11332, A2 => n11565, B1 => n8508, B2 => 
                           n11452, ZN => n2067);
   U10151 : OAI22_X1 port map( A1 => n11332, A2 => n11569, B1 => n8507, B2 => 
                           n11452, ZN => n2068);
   U10152 : OAI22_X1 port map( A1 => n11332, A2 => n11573, B1 => n8506, B2 => 
                           n11452, ZN => n2069);
   U10153 : OAI22_X1 port map( A1 => n11332, A2 => n11577, B1 => n8505, B2 => 
                           n10524, ZN => n2070);
   U10154 : OAI22_X1 port map( A1 => n11332, A2 => n11581, B1 => n8504, B2 => 
                           n10524, ZN => n2071);
   U10155 : OAI22_X1 port map( A1 => n11332, A2 => n11585, B1 => n8503, B2 => 
                           n10524, ZN => n2072);
   U10156 : OAI22_X1 port map( A1 => n11332, A2 => n11589, B1 => n8502, B2 => 
                           n10524, ZN => n2073);
   U10157 : OAI22_X1 port map( A1 => n11332, A2 => n11593, B1 => n8501, B2 => 
                           n10524, ZN => n2074);
   U10158 : OAI22_X1 port map( A1 => n11332, A2 => n11597, B1 => n8500, B2 => 
                           n10524, ZN => n2075);
   U10159 : OAI22_X1 port map( A1 => n11332, A2 => n11601, B1 => n8499, B2 => 
                           n10524, ZN => n2076);
   U10160 : OAI22_X1 port map( A1 => n11332, A2 => n11609, B1 => n8498, B2 => 
                           n10524, ZN => n2077);
   U10161 : OAI22_X1 port map( A1 => n11346, A2 => n11481, B1 => n8401, B2 => 
                           n11468, ZN => n2174);
   U10162 : OAI22_X1 port map( A1 => n11346, A2 => n11485, B1 => n8400, B2 => 
                           n11468, ZN => n2175);
   U10163 : OAI22_X1 port map( A1 => n11346, A2 => n11489, B1 => n8399, B2 => 
                           n11468, ZN => n2176);
   U10164 : OAI22_X1 port map( A1 => n11346, A2 => n11493, B1 => n8398, B2 => 
                           n11468, ZN => n2177);
   U10165 : OAI22_X1 port map( A1 => n11346, A2 => n11497, B1 => n8397, B2 => 
                           n11468, ZN => n2178);
   U10166 : OAI22_X1 port map( A1 => n11346, A2 => n11501, B1 => n8396, B2 => 
                           n11468, ZN => n2179);
   U10167 : OAI22_X1 port map( A1 => n11346, A2 => n11505, B1 => n8395, B2 => 
                           n11468, ZN => n2180);
   U10168 : OAI22_X1 port map( A1 => n11346, A2 => n11509, B1 => n8394, B2 => 
                           n11468, ZN => n2181);
   U10169 : OAI22_X1 port map( A1 => n11345, A2 => n11513, B1 => n8393, B2 => 
                           n11468, ZN => n2182);
   U10170 : OAI22_X1 port map( A1 => n11345, A2 => n11517, B1 => n8392, B2 => 
                           n11468, ZN => n2183);
   U10171 : OAI22_X1 port map( A1 => n11345, A2 => n11521, B1 => n8391, B2 => 
                           n11468, ZN => n2184);
   U10172 : OAI22_X1 port map( A1 => n11345, A2 => n11525, B1 => n8390, B2 => 
                           n11468, ZN => n2185);
   U10173 : OAI22_X1 port map( A1 => n11345, A2 => n11529, B1 => n8389, B2 => 
                           n10517, ZN => n2186);
   U10174 : OAI22_X1 port map( A1 => n11345, A2 => n11533, B1 => n8388, B2 => 
                           n10517, ZN => n2187);
   U10175 : OAI22_X1 port map( A1 => n11345, A2 => n11537, B1 => n8387, B2 => 
                           n10517, ZN => n2188);
   U10176 : OAI22_X1 port map( A1 => n11345, A2 => n11541, B1 => n8386, B2 => 
                           n11468, ZN => n2189);
   U10177 : OAI22_X1 port map( A1 => n11345, A2 => n11545, B1 => n8385, B2 => 
                           n11468, ZN => n2190);
   U10178 : OAI22_X1 port map( A1 => n11345, A2 => n11549, B1 => n8384, B2 => 
                           n11468, ZN => n2191);
   U10179 : OAI22_X1 port map( A1 => n11345, A2 => n11553, B1 => n8383, B2 => 
                           n11468, ZN => n2192);
   U10180 : OAI22_X1 port map( A1 => n11345, A2 => n11557, B1 => n8382, B2 => 
                           n11468, ZN => n2193);
   U10181 : OAI22_X1 port map( A1 => n11344, A2 => n11561, B1 => n8381, B2 => 
                           n11468, ZN => n2194);
   U10182 : OAI22_X1 port map( A1 => n11344, A2 => n11565, B1 => n8380, B2 => 
                           n11468, ZN => n2195);
   U10183 : OAI22_X1 port map( A1 => n11344, A2 => n11569, B1 => n8379, B2 => 
                           n11468, ZN => n2196);
   U10184 : OAI22_X1 port map( A1 => n11344, A2 => n11573, B1 => n8378, B2 => 
                           n11468, ZN => n2197);
   U10185 : OAI22_X1 port map( A1 => n11344, A2 => n11577, B1 => n8377, B2 => 
                           n10517, ZN => n2198);
   U10186 : OAI22_X1 port map( A1 => n11344, A2 => n11581, B1 => n8376, B2 => 
                           n10517, ZN => n2199);
   U10187 : OAI22_X1 port map( A1 => n11344, A2 => n11585, B1 => n8375, B2 => 
                           n10517, ZN => n2200);
   U10188 : OAI22_X1 port map( A1 => n11344, A2 => n11589, B1 => n8374, B2 => 
                           n10517, ZN => n2201);
   U10189 : OAI22_X1 port map( A1 => n11344, A2 => n11593, B1 => n8373, B2 => 
                           n10517, ZN => n2202);
   U10190 : OAI22_X1 port map( A1 => n11344, A2 => n11597, B1 => n8372, B2 => 
                           n10517, ZN => n2203);
   U10191 : OAI22_X1 port map( A1 => n11344, A2 => n11601, B1 => n8371, B2 => 
                           n10517, ZN => n2204);
   U10192 : OAI22_X1 port map( A1 => n11344, A2 => n11609, B1 => n8370, B2 => 
                           n10517, ZN => n2205);
   U10193 : OAI22_X1 port map( A1 => n11277, A2 => n11483, B1 => n9137, B2 => 
                           n11376, ZN => n1438);
   U10194 : OAI22_X1 port map( A1 => n11277, A2 => n11487, B1 => n9136, B2 => 
                           n11376, ZN => n1439);
   U10195 : OAI22_X1 port map( A1 => n11277, A2 => n11491, B1 => n9135, B2 => 
                           n11376, ZN => n1440);
   U10196 : OAI22_X1 port map( A1 => n11277, A2 => n11495, B1 => n9134, B2 => 
                           n11376, ZN => n1441);
   U10197 : OAI22_X1 port map( A1 => n11277, A2 => n11499, B1 => n9133, B2 => 
                           n11376, ZN => n1442);
   U10198 : OAI22_X1 port map( A1 => n11277, A2 => n11503, B1 => n9132, B2 => 
                           n11376, ZN => n1443);
   U10199 : OAI22_X1 port map( A1 => n11277, A2 => n11507, B1 => n9131, B2 => 
                           n11376, ZN => n1444);
   U10200 : OAI22_X1 port map( A1 => n11277, A2 => n11511, B1 => n9130, B2 => 
                           n11376, ZN => n1445);
   U10201 : OAI22_X1 port map( A1 => n11276, A2 => n11515, B1 => n9129, B2 => 
                           n11376, ZN => n1446);
   U10202 : OAI22_X1 port map( A1 => n11276, A2 => n11519, B1 => n9128, B2 => 
                           n11376, ZN => n1447);
   U10203 : OAI22_X1 port map( A1 => n11276, A2 => n11523, B1 => n9127, B2 => 
                           n11376, ZN => n1448);
   U10204 : OAI22_X1 port map( A1 => n11276, A2 => n11527, B1 => n9126, B2 => 
                           n11376, ZN => n1449);
   U10205 : OAI22_X1 port map( A1 => n11276, A2 => n11531, B1 => n9125, B2 => 
                           n10549, ZN => n1450);
   U10206 : OAI22_X1 port map( A1 => n11276, A2 => n11535, B1 => n9124, B2 => 
                           n10549, ZN => n1451);
   U10207 : OAI22_X1 port map( A1 => n11276, A2 => n11539, B1 => n9123, B2 => 
                           n10549, ZN => n1452);
   U10208 : OAI22_X1 port map( A1 => n11276, A2 => n11543, B1 => n9122, B2 => 
                           n11376, ZN => n1453);
   U10209 : OAI22_X1 port map( A1 => n11276, A2 => n11547, B1 => n9121, B2 => 
                           n11376, ZN => n1454);
   U10210 : OAI22_X1 port map( A1 => n11276, A2 => n11551, B1 => n9120, B2 => 
                           n11376, ZN => n1455);
   U10211 : OAI22_X1 port map( A1 => n11276, A2 => n11555, B1 => n9119, B2 => 
                           n11376, ZN => n1456);
   U10212 : OAI22_X1 port map( A1 => n11276, A2 => n11559, B1 => n9118, B2 => 
                           n11376, ZN => n1457);
   U10213 : OAI22_X1 port map( A1 => n11275, A2 => n11563, B1 => n9117, B2 => 
                           n11376, ZN => n1458);
   U10214 : OAI22_X1 port map( A1 => n11275, A2 => n11567, B1 => n9116, B2 => 
                           n11376, ZN => n1459);
   U10215 : OAI22_X1 port map( A1 => n11275, A2 => n11571, B1 => n9115, B2 => 
                           n11376, ZN => n1460);
   U10216 : OAI22_X1 port map( A1 => n11275, A2 => n11575, B1 => n9114, B2 => 
                           n11376, ZN => n1461);
   U10217 : OAI22_X1 port map( A1 => n11275, A2 => n11579, B1 => n9113, B2 => 
                           n10549, ZN => n1462);
   U10218 : OAI22_X1 port map( A1 => n11275, A2 => n11583, B1 => n9112, B2 => 
                           n10549, ZN => n1463);
   U10219 : OAI22_X1 port map( A1 => n11275, A2 => n11587, B1 => n9111, B2 => 
                           n10549, ZN => n1464);
   U10220 : OAI22_X1 port map( A1 => n11275, A2 => n11591, B1 => n9110, B2 => 
                           n10549, ZN => n1465);
   U10221 : OAI22_X1 port map( A1 => n11275, A2 => n11595, B1 => n9109, B2 => 
                           n10549, ZN => n1466);
   U10222 : OAI22_X1 port map( A1 => n11275, A2 => n11599, B1 => n9108, B2 => 
                           n10549, ZN => n1467);
   U10223 : OAI22_X1 port map( A1 => n11275, A2 => n11603, B1 => n9107, B2 => 
                           n10549, ZN => n1468);
   U10224 : OAI22_X1 port map( A1 => n11275, A2 => n11611, B1 => n9106, B2 => 
                           n10549, ZN => n1469);
   U10225 : OAI22_X1 port map( A1 => n11289, A2 => n11482, B1 => n9009, B2 => 
                           n11392, ZN => n1566);
   U10226 : OAI22_X1 port map( A1 => n11289, A2 => n11486, B1 => n9008, B2 => 
                           n11392, ZN => n1567);
   U10227 : OAI22_X1 port map( A1 => n11289, A2 => n11490, B1 => n9007, B2 => 
                           n11392, ZN => n1568);
   U10228 : OAI22_X1 port map( A1 => n11289, A2 => n11494, B1 => n9006, B2 => 
                           n11392, ZN => n1569);
   U10229 : OAI22_X1 port map( A1 => n11289, A2 => n11498, B1 => n9005, B2 => 
                           n11392, ZN => n1570);
   U10230 : OAI22_X1 port map( A1 => n11289, A2 => n11502, B1 => n9004, B2 => 
                           n11392, ZN => n1571);
   U10231 : OAI22_X1 port map( A1 => n11289, A2 => n11506, B1 => n9003, B2 => 
                           n11392, ZN => n1572);
   U10232 : OAI22_X1 port map( A1 => n11289, A2 => n11510, B1 => n9002, B2 => 
                           n11392, ZN => n1573);
   U10233 : OAI22_X1 port map( A1 => n11288, A2 => n11514, B1 => n9001, B2 => 
                           n11392, ZN => n1574);
   U10234 : OAI22_X1 port map( A1 => n11288, A2 => n11518, B1 => n9000, B2 => 
                           n11392, ZN => n1575);
   U10235 : OAI22_X1 port map( A1 => n11288, A2 => n11522, B1 => n8999, B2 => 
                           n11392, ZN => n1576);
   U10236 : OAI22_X1 port map( A1 => n11288, A2 => n11526, B1 => n8998, B2 => 
                           n11392, ZN => n1577);
   U10237 : OAI22_X1 port map( A1 => n11288, A2 => n11530, B1 => n8997, B2 => 
                           n10544, ZN => n1578);
   U10238 : OAI22_X1 port map( A1 => n11288, A2 => n11534, B1 => n8996, B2 => 
                           n10544, ZN => n1579);
   U10239 : OAI22_X1 port map( A1 => n11288, A2 => n11538, B1 => n8995, B2 => 
                           n10544, ZN => n1580);
   U10240 : OAI22_X1 port map( A1 => n11288, A2 => n11542, B1 => n8994, B2 => 
                           n11392, ZN => n1581);
   U10241 : OAI22_X1 port map( A1 => n11288, A2 => n11546, B1 => n8993, B2 => 
                           n11392, ZN => n1582);
   U10242 : OAI22_X1 port map( A1 => n11288, A2 => n11550, B1 => n8992, B2 => 
                           n11392, ZN => n1583);
   U10243 : OAI22_X1 port map( A1 => n11288, A2 => n11554, B1 => n8991, B2 => 
                           n11392, ZN => n1584);
   U10244 : OAI22_X1 port map( A1 => n11288, A2 => n11558, B1 => n8990, B2 => 
                           n11392, ZN => n1585);
   U10245 : OAI22_X1 port map( A1 => n11287, A2 => n11562, B1 => n8989, B2 => 
                           n11392, ZN => n1586);
   U10246 : OAI22_X1 port map( A1 => n11287, A2 => n11566, B1 => n8988, B2 => 
                           n11392, ZN => n1587);
   U10247 : OAI22_X1 port map( A1 => n11287, A2 => n11570, B1 => n8987, B2 => 
                           n11392, ZN => n1588);
   U10248 : OAI22_X1 port map( A1 => n11287, A2 => n11574, B1 => n8986, B2 => 
                           n11392, ZN => n1589);
   U10249 : OAI22_X1 port map( A1 => n11287, A2 => n11578, B1 => n8985, B2 => 
                           n10544, ZN => n1590);
   U10250 : OAI22_X1 port map( A1 => n11287, A2 => n11582, B1 => n8984, B2 => 
                           n10544, ZN => n1591);
   U10251 : OAI22_X1 port map( A1 => n11287, A2 => n11586, B1 => n8983, B2 => 
                           n10544, ZN => n1592);
   U10252 : OAI22_X1 port map( A1 => n11287, A2 => n11590, B1 => n8982, B2 => 
                           n10544, ZN => n1593);
   U10253 : OAI22_X1 port map( A1 => n11287, A2 => n11594, B1 => n8981, B2 => 
                           n10544, ZN => n1594);
   U10254 : OAI22_X1 port map( A1 => n11287, A2 => n11598, B1 => n8980, B2 => 
                           n10544, ZN => n1595);
   U10255 : OAI22_X1 port map( A1 => n11287, A2 => n11602, B1 => n8979, B2 => 
                           n10544, ZN => n1596);
   U10256 : OAI22_X1 port map( A1 => n11287, A2 => n11610, B1 => n8978, B2 => 
                           n10544, ZN => n1597);
   U10257 : OAI22_X1 port map( A1 => n11304, A2 => n11482, B1 => n8849, B2 => 
                           n11412, ZN => n1726);
   U10258 : OAI22_X1 port map( A1 => n11304, A2 => n11486, B1 => n8848, B2 => 
                           n11412, ZN => n1727);
   U10259 : OAI22_X1 port map( A1 => n11304, A2 => n11490, B1 => n8847, B2 => 
                           n11412, ZN => n1728);
   U10260 : OAI22_X1 port map( A1 => n11304, A2 => n11494, B1 => n8846, B2 => 
                           n11412, ZN => n1729);
   U10261 : OAI22_X1 port map( A1 => n11304, A2 => n11498, B1 => n8845, B2 => 
                           n11412, ZN => n1730);
   U10262 : OAI22_X1 port map( A1 => n11304, A2 => n11502, B1 => n8844, B2 => 
                           n11412, ZN => n1731);
   U10263 : OAI22_X1 port map( A1 => n11304, A2 => n11506, B1 => n8843, B2 => 
                           n11412, ZN => n1732);
   U10264 : OAI22_X1 port map( A1 => n11304, A2 => n11510, B1 => n8842, B2 => 
                           n11412, ZN => n1733);
   U10265 : OAI22_X1 port map( A1 => n11303, A2 => n11514, B1 => n8841, B2 => 
                           n11412, ZN => n1734);
   U10266 : OAI22_X1 port map( A1 => n11303, A2 => n11518, B1 => n8840, B2 => 
                           n11412, ZN => n1735);
   U10267 : OAI22_X1 port map( A1 => n11303, A2 => n11522, B1 => n8839, B2 => 
                           n11412, ZN => n1736);
   U10268 : OAI22_X1 port map( A1 => n11303, A2 => n11526, B1 => n8838, B2 => 
                           n11412, ZN => n1737);
   U10269 : OAI22_X1 port map( A1 => n11303, A2 => n11530, B1 => n8837, B2 => 
                           n10537, ZN => n1738);
   U10270 : OAI22_X1 port map( A1 => n11303, A2 => n11534, B1 => n8836, B2 => 
                           n10537, ZN => n1739);
   U10271 : OAI22_X1 port map( A1 => n11303, A2 => n11538, B1 => n8835, B2 => 
                           n10537, ZN => n1740);
   U10272 : OAI22_X1 port map( A1 => n11303, A2 => n11542, B1 => n8834, B2 => 
                           n11412, ZN => n1741);
   U10273 : OAI22_X1 port map( A1 => n11303, A2 => n11546, B1 => n8833, B2 => 
                           n11412, ZN => n1742);
   U10274 : OAI22_X1 port map( A1 => n11303, A2 => n11550, B1 => n8832, B2 => 
                           n11412, ZN => n1743);
   U10275 : OAI22_X1 port map( A1 => n11303, A2 => n11554, B1 => n8831, B2 => 
                           n11412, ZN => n1744);
   U10276 : OAI22_X1 port map( A1 => n11303, A2 => n11558, B1 => n8830, B2 => 
                           n11412, ZN => n1745);
   U10277 : OAI22_X1 port map( A1 => n11302, A2 => n11562, B1 => n8829, B2 => 
                           n11412, ZN => n1746);
   U10278 : OAI22_X1 port map( A1 => n11302, A2 => n11566, B1 => n8828, B2 => 
                           n11412, ZN => n1747);
   U10279 : OAI22_X1 port map( A1 => n11302, A2 => n11570, B1 => n8827, B2 => 
                           n11412, ZN => n1748);
   U10280 : OAI22_X1 port map( A1 => n11302, A2 => n11574, B1 => n8826, B2 => 
                           n11412, ZN => n1749);
   U10281 : OAI22_X1 port map( A1 => n11302, A2 => n11578, B1 => n8825, B2 => 
                           n10537, ZN => n1750);
   U10282 : OAI22_X1 port map( A1 => n11302, A2 => n11582, B1 => n8824, B2 => 
                           n10537, ZN => n1751);
   U10283 : OAI22_X1 port map( A1 => n11302, A2 => n11586, B1 => n8823, B2 => 
                           n10537, ZN => n1752);
   U10284 : OAI22_X1 port map( A1 => n11302, A2 => n11590, B1 => n8822, B2 => 
                           n10537, ZN => n1753);
   U10285 : OAI22_X1 port map( A1 => n11302, A2 => n11594, B1 => n8821, B2 => 
                           n10537, ZN => n1754);
   U10286 : OAI22_X1 port map( A1 => n11302, A2 => n11598, B1 => n8820, B2 => 
                           n10537, ZN => n1755);
   U10287 : OAI22_X1 port map( A1 => n11302, A2 => n11602, B1 => n8819, B2 => 
                           n10537, ZN => n1756);
   U10288 : OAI22_X1 port map( A1 => n11302, A2 => n11610, B1 => n8818, B2 => 
                           n10537, ZN => n1757);
   U10289 : OAI22_X1 port map( A1 => n11310, A2 => n11482, B1 => n8785, B2 => 
                           n11420, ZN => n1790);
   U10290 : OAI22_X1 port map( A1 => n11310, A2 => n11486, B1 => n8784, B2 => 
                           n11420, ZN => n1791);
   U10291 : OAI22_X1 port map( A1 => n11310, A2 => n11490, B1 => n8783, B2 => 
                           n11420, ZN => n1792);
   U10292 : OAI22_X1 port map( A1 => n11310, A2 => n11494, B1 => n8782, B2 => 
                           n11420, ZN => n1793);
   U10293 : OAI22_X1 port map( A1 => n11310, A2 => n11498, B1 => n8781, B2 => 
                           n11420, ZN => n1794);
   U10294 : OAI22_X1 port map( A1 => n11310, A2 => n11502, B1 => n8780, B2 => 
                           n11420, ZN => n1795);
   U10295 : OAI22_X1 port map( A1 => n11310, A2 => n11506, B1 => n8779, B2 => 
                           n11420, ZN => n1796);
   U10296 : OAI22_X1 port map( A1 => n11310, A2 => n11510, B1 => n8778, B2 => 
                           n11420, ZN => n1797);
   U10297 : OAI22_X1 port map( A1 => n11309, A2 => n11514, B1 => n8777, B2 => 
                           n11420, ZN => n1798);
   U10298 : OAI22_X1 port map( A1 => n11309, A2 => n11518, B1 => n8776, B2 => 
                           n11420, ZN => n1799);
   U10299 : OAI22_X1 port map( A1 => n11309, A2 => n11522, B1 => n8775, B2 => 
                           n11420, ZN => n1800);
   U10300 : OAI22_X1 port map( A1 => n11309, A2 => n11526, B1 => n8774, B2 => 
                           n11420, ZN => n1801);
   U10301 : OAI22_X1 port map( A1 => n11309, A2 => n11530, B1 => n8773, B2 => 
                           n10534, ZN => n1802);
   U10302 : OAI22_X1 port map( A1 => n11309, A2 => n11534, B1 => n8772, B2 => 
                           n10534, ZN => n1803);
   U10303 : OAI22_X1 port map( A1 => n11309, A2 => n11538, B1 => n8771, B2 => 
                           n10534, ZN => n1804);
   U10304 : OAI22_X1 port map( A1 => n11309, A2 => n11542, B1 => n8770, B2 => 
                           n11420, ZN => n1805);
   U10305 : OAI22_X1 port map( A1 => n11309, A2 => n11546, B1 => n8769, B2 => 
                           n11420, ZN => n1806);
   U10306 : OAI22_X1 port map( A1 => n11309, A2 => n11550, B1 => n8768, B2 => 
                           n11420, ZN => n1807);
   U10307 : OAI22_X1 port map( A1 => n11309, A2 => n11554, B1 => n8767, B2 => 
                           n11420, ZN => n1808);
   U10308 : OAI22_X1 port map( A1 => n11309, A2 => n11558, B1 => n8766, B2 => 
                           n11420, ZN => n1809);
   U10309 : OAI22_X1 port map( A1 => n11308, A2 => n11562, B1 => n8765, B2 => 
                           n11420, ZN => n1810);
   U10310 : OAI22_X1 port map( A1 => n11308, A2 => n11566, B1 => n8764, B2 => 
                           n11420, ZN => n1811);
   U10311 : OAI22_X1 port map( A1 => n11308, A2 => n11570, B1 => n8763, B2 => 
                           n11420, ZN => n1812);
   U10312 : OAI22_X1 port map( A1 => n11308, A2 => n11574, B1 => n8762, B2 => 
                           n11420, ZN => n1813);
   U10313 : OAI22_X1 port map( A1 => n11308, A2 => n11578, B1 => n8761, B2 => 
                           n10534, ZN => n1814);
   U10314 : OAI22_X1 port map( A1 => n11308, A2 => n11582, B1 => n8760, B2 => 
                           n10534, ZN => n1815);
   U10315 : OAI22_X1 port map( A1 => n11308, A2 => n11586, B1 => n8759, B2 => 
                           n10534, ZN => n1816);
   U10316 : OAI22_X1 port map( A1 => n11308, A2 => n11590, B1 => n8758, B2 => 
                           n10534, ZN => n1817);
   U10317 : OAI22_X1 port map( A1 => n11308, A2 => n11594, B1 => n8757, B2 => 
                           n10534, ZN => n1818);
   U10318 : OAI22_X1 port map( A1 => n11308, A2 => n11598, B1 => n8756, B2 => 
                           n10534, ZN => n1819);
   U10319 : OAI22_X1 port map( A1 => n11308, A2 => n11602, B1 => n8755, B2 => 
                           n10534, ZN => n1820);
   U10320 : OAI22_X1 port map( A1 => n11308, A2 => n11610, B1 => n8754, B2 => 
                           n10534, ZN => n1821);
   U10321 : OAI22_X1 port map( A1 => n11328, A2 => n11481, B1 => n8593, B2 => 
                           n11444, ZN => n1982);
   U10322 : OAI22_X1 port map( A1 => n11328, A2 => n11485, B1 => n8592, B2 => 
                           n11444, ZN => n1983);
   U10323 : OAI22_X1 port map( A1 => n11328, A2 => n11489, B1 => n8591, B2 => 
                           n11444, ZN => n1984);
   U10324 : OAI22_X1 port map( A1 => n11328, A2 => n11493, B1 => n8590, B2 => 
                           n11444, ZN => n1985);
   U10325 : OAI22_X1 port map( A1 => n11328, A2 => n11497, B1 => n8589, B2 => 
                           n11444, ZN => n1986);
   U10326 : OAI22_X1 port map( A1 => n11328, A2 => n11501, B1 => n8588, B2 => 
                           n11444, ZN => n1987);
   U10327 : OAI22_X1 port map( A1 => n11328, A2 => n11505, B1 => n8587, B2 => 
                           n11444, ZN => n1988);
   U10328 : OAI22_X1 port map( A1 => n11328, A2 => n11509, B1 => n8586, B2 => 
                           n11444, ZN => n1989);
   U10329 : OAI22_X1 port map( A1 => n11327, A2 => n11513, B1 => n8585, B2 => 
                           n11444, ZN => n1990);
   U10330 : OAI22_X1 port map( A1 => n11327, A2 => n11517, B1 => n8584, B2 => 
                           n11444, ZN => n1991);
   U10331 : OAI22_X1 port map( A1 => n11327, A2 => n11521, B1 => n8583, B2 => 
                           n11444, ZN => n1992);
   U10332 : OAI22_X1 port map( A1 => n11327, A2 => n11525, B1 => n8582, B2 => 
                           n11444, ZN => n1993);
   U10333 : OAI22_X1 port map( A1 => n11327, A2 => n11529, B1 => n8581, B2 => 
                           n10527, ZN => n1994);
   U10334 : OAI22_X1 port map( A1 => n11327, A2 => n11533, B1 => n8580, B2 => 
                           n10527, ZN => n1995);
   U10335 : OAI22_X1 port map( A1 => n11327, A2 => n11537, B1 => n8579, B2 => 
                           n10527, ZN => n1996);
   U10336 : OAI22_X1 port map( A1 => n11327, A2 => n11541, B1 => n8578, B2 => 
                           n11444, ZN => n1997);
   U10337 : OAI22_X1 port map( A1 => n11327, A2 => n11545, B1 => n8577, B2 => 
                           n11444, ZN => n1998);
   U10338 : OAI22_X1 port map( A1 => n11327, A2 => n11549, B1 => n8576, B2 => 
                           n11444, ZN => n1999);
   U10339 : OAI22_X1 port map( A1 => n11327, A2 => n11553, B1 => n8575, B2 => 
                           n11444, ZN => n2000);
   U10340 : OAI22_X1 port map( A1 => n11327, A2 => n11557, B1 => n8574, B2 => 
                           n11444, ZN => n2001);
   U10341 : OAI22_X1 port map( A1 => n11326, A2 => n11561, B1 => n8573, B2 => 
                           n11444, ZN => n2002);
   U10342 : OAI22_X1 port map( A1 => n11326, A2 => n11565, B1 => n8572, B2 => 
                           n11444, ZN => n2003);
   U10343 : OAI22_X1 port map( A1 => n11326, A2 => n11569, B1 => n8571, B2 => 
                           n11444, ZN => n2004);
   U10344 : OAI22_X1 port map( A1 => n11326, A2 => n11573, B1 => n8570, B2 => 
                           n11444, ZN => n2005);
   U10345 : OAI22_X1 port map( A1 => n11326, A2 => n11577, B1 => n8569, B2 => 
                           n10527, ZN => n2006);
   U10346 : OAI22_X1 port map( A1 => n11326, A2 => n11581, B1 => n8568, B2 => 
                           n10527, ZN => n2007);
   U10347 : OAI22_X1 port map( A1 => n11326, A2 => n11585, B1 => n8567, B2 => 
                           n10527, ZN => n2008);
   U10348 : OAI22_X1 port map( A1 => n11326, A2 => n11589, B1 => n8566, B2 => 
                           n10527, ZN => n2009);
   U10349 : OAI22_X1 port map( A1 => n11326, A2 => n11593, B1 => n8565, B2 => 
                           n10527, ZN => n2010);
   U10350 : OAI22_X1 port map( A1 => n11326, A2 => n11597, B1 => n8564, B2 => 
                           n10527, ZN => n2011);
   U10351 : OAI22_X1 port map( A1 => n11326, A2 => n11601, B1 => n8563, B2 => 
                           n10527, ZN => n2012);
   U10352 : OAI22_X1 port map( A1 => n11326, A2 => n11609, B1 => n8562, B2 => 
                           n10527, ZN => n2013);
   U10353 : OAI22_X1 port map( A1 => n11337, A2 => n11481, B1 => n8497, B2 => 
                           n11456, ZN => n2078);
   U10354 : OAI22_X1 port map( A1 => n11337, A2 => n11485, B1 => n8496, B2 => 
                           n11456, ZN => n2079);
   U10355 : OAI22_X1 port map( A1 => n11337, A2 => n11489, B1 => n8495, B2 => 
                           n11456, ZN => n2080);
   U10356 : OAI22_X1 port map( A1 => n11337, A2 => n11493, B1 => n8494, B2 => 
                           n11456, ZN => n2081);
   U10357 : OAI22_X1 port map( A1 => n11337, A2 => n11497, B1 => n8493, B2 => 
                           n11456, ZN => n2082);
   U10358 : OAI22_X1 port map( A1 => n11337, A2 => n11501, B1 => n8492, B2 => 
                           n11456, ZN => n2083);
   U10359 : OAI22_X1 port map( A1 => n11337, A2 => n11505, B1 => n8491, B2 => 
                           n11456, ZN => n2084);
   U10360 : OAI22_X1 port map( A1 => n11337, A2 => n11509, B1 => n8490, B2 => 
                           n11456, ZN => n2085);
   U10361 : OAI22_X1 port map( A1 => n11336, A2 => n11513, B1 => n8489, B2 => 
                           n11456, ZN => n2086);
   U10362 : OAI22_X1 port map( A1 => n11336, A2 => n11517, B1 => n8488, B2 => 
                           n11456, ZN => n2087);
   U10363 : OAI22_X1 port map( A1 => n11336, A2 => n11521, B1 => n8487, B2 => 
                           n11456, ZN => n2088);
   U10364 : OAI22_X1 port map( A1 => n11336, A2 => n11525, B1 => n8486, B2 => 
                           n11456, ZN => n2089);
   U10365 : OAI22_X1 port map( A1 => n11336, A2 => n11529, B1 => n8485, B2 => 
                           n10523, ZN => n2090);
   U10366 : OAI22_X1 port map( A1 => n11336, A2 => n11533, B1 => n8484, B2 => 
                           n10523, ZN => n2091);
   U10367 : OAI22_X1 port map( A1 => n11336, A2 => n11537, B1 => n8483, B2 => 
                           n10523, ZN => n2092);
   U10368 : OAI22_X1 port map( A1 => n11336, A2 => n11541, B1 => n8482, B2 => 
                           n11456, ZN => n2093);
   U10369 : OAI22_X1 port map( A1 => n11336, A2 => n11545, B1 => n8481, B2 => 
                           n11456, ZN => n2094);
   U10370 : OAI22_X1 port map( A1 => n11336, A2 => n11549, B1 => n8480, B2 => 
                           n11456, ZN => n2095);
   U10371 : OAI22_X1 port map( A1 => n11336, A2 => n11553, B1 => n8479, B2 => 
                           n11456, ZN => n2096);
   U10372 : OAI22_X1 port map( A1 => n11336, A2 => n11557, B1 => n8478, B2 => 
                           n11456, ZN => n2097);
   U10373 : OAI22_X1 port map( A1 => n11335, A2 => n11561, B1 => n8477, B2 => 
                           n11456, ZN => n2098);
   U10374 : OAI22_X1 port map( A1 => n11335, A2 => n11565, B1 => n8476, B2 => 
                           n11456, ZN => n2099);
   U10375 : OAI22_X1 port map( A1 => n11335, A2 => n11569, B1 => n8475, B2 => 
                           n11456, ZN => n2100);
   U10376 : OAI22_X1 port map( A1 => n11335, A2 => n11573, B1 => n8474, B2 => 
                           n11456, ZN => n2101);
   U10377 : OAI22_X1 port map( A1 => n11335, A2 => n11577, B1 => n8473, B2 => 
                           n10523, ZN => n2102);
   U10378 : OAI22_X1 port map( A1 => n11335, A2 => n11581, B1 => n8472, B2 => 
                           n10523, ZN => n2103);
   U10379 : OAI22_X1 port map( A1 => n11335, A2 => n11585, B1 => n8471, B2 => 
                           n10523, ZN => n2104);
   U10380 : OAI22_X1 port map( A1 => n11335, A2 => n11589, B1 => n8470, B2 => 
                           n10523, ZN => n2105);
   U10381 : OAI22_X1 port map( A1 => n11335, A2 => n11593, B1 => n8469, B2 => 
                           n10523, ZN => n2106);
   U10382 : OAI22_X1 port map( A1 => n11335, A2 => n11597, B1 => n8468, B2 => 
                           n10523, ZN => n2107);
   U10383 : OAI22_X1 port map( A1 => n11335, A2 => n11601, B1 => n8467, B2 => 
                           n10523, ZN => n2108);
   U10384 : OAI22_X1 port map( A1 => n11335, A2 => n11609, B1 => n8466, B2 => 
                           n10523, ZN => n2109);
   U10385 : OAI22_X1 port map( A1 => n11355, A2 => n11481, B1 => n8305, B2 => 
                           n11604, ZN => n2270);
   U10386 : OAI22_X1 port map( A1 => n11355, A2 => n11485, B1 => n8304, B2 => 
                           n11604, ZN => n2271);
   U10387 : OAI22_X1 port map( A1 => n11355, A2 => n11489, B1 => n8303, B2 => 
                           n11604, ZN => n2272);
   U10388 : OAI22_X1 port map( A1 => n11355, A2 => n11493, B1 => n8302, B2 => 
                           n11604, ZN => n2273);
   U10389 : OAI22_X1 port map( A1 => n11355, A2 => n11497, B1 => n8301, B2 => 
                           n11604, ZN => n2274);
   U10390 : OAI22_X1 port map( A1 => n11355, A2 => n11501, B1 => n8300, B2 => 
                           n11604, ZN => n2275);
   U10391 : OAI22_X1 port map( A1 => n11355, A2 => n11505, B1 => n8299, B2 => 
                           n11604, ZN => n2276);
   U10392 : OAI22_X1 port map( A1 => n11355, A2 => n11509, B1 => n8298, B2 => 
                           n11604, ZN => n2277);
   U10393 : OAI22_X1 port map( A1 => n11354, A2 => n11513, B1 => n8297, B2 => 
                           n11604, ZN => n2278);
   U10394 : OAI22_X1 port map( A1 => n11354, A2 => n11517, B1 => n8296, B2 => 
                           n11604, ZN => n2279);
   U10395 : OAI22_X1 port map( A1 => n11354, A2 => n11521, B1 => n8295, B2 => 
                           n11604, ZN => n2280);
   U10396 : OAI22_X1 port map( A1 => n11354, A2 => n11525, B1 => n8294, B2 => 
                           n11604, ZN => n2281);
   U10397 : OAI22_X1 port map( A1 => n11354, A2 => n11529, B1 => n8293, B2 => 
                           n10479, ZN => n2282);
   U10398 : OAI22_X1 port map( A1 => n11354, A2 => n11533, B1 => n8292, B2 => 
                           n10479, ZN => n2283);
   U10399 : OAI22_X1 port map( A1 => n11354, A2 => n11537, B1 => n8291, B2 => 
                           n10479, ZN => n2284);
   U10400 : OAI22_X1 port map( A1 => n11354, A2 => n11541, B1 => n8290, B2 => 
                           n11604, ZN => n2285);
   U10401 : OAI22_X1 port map( A1 => n11354, A2 => n11545, B1 => n8289, B2 => 
                           n11604, ZN => n2286);
   U10402 : OAI22_X1 port map( A1 => n11354, A2 => n11549, B1 => n8288, B2 => 
                           n11604, ZN => n2287);
   U10403 : OAI22_X1 port map( A1 => n11354, A2 => n11553, B1 => n8287, B2 => 
                           n11604, ZN => n2288);
   U10404 : OAI22_X1 port map( A1 => n11354, A2 => n11557, B1 => n8286, B2 => 
                           n11604, ZN => n2289);
   U10405 : OAI22_X1 port map( A1 => n11353, A2 => n11561, B1 => n8285, B2 => 
                           n11604, ZN => n2290);
   U10406 : OAI22_X1 port map( A1 => n11353, A2 => n11565, B1 => n8284, B2 => 
                           n11604, ZN => n2291);
   U10407 : OAI22_X1 port map( A1 => n11353, A2 => n11569, B1 => n8283, B2 => 
                           n11604, ZN => n2292);
   U10408 : OAI22_X1 port map( A1 => n11353, A2 => n11573, B1 => n8282, B2 => 
                           n11604, ZN => n2293);
   U10409 : OAI22_X1 port map( A1 => n11353, A2 => n11577, B1 => n8281, B2 => 
                           n10479, ZN => n2294);
   U10410 : OAI22_X1 port map( A1 => n11353, A2 => n11581, B1 => n8280, B2 => 
                           n10479, ZN => n2295);
   U10411 : OAI22_X1 port map( A1 => n11353, A2 => n11585, B1 => n8279, B2 => 
                           n10479, ZN => n2296);
   U10412 : OAI22_X1 port map( A1 => n11353, A2 => n11589, B1 => n8278, B2 => 
                           n10479, ZN => n2297);
   U10413 : OAI22_X1 port map( A1 => n11353, A2 => n11593, B1 => n8277, B2 => 
                           n10479, ZN => n2298);
   U10414 : OAI22_X1 port map( A1 => n11353, A2 => n11597, B1 => n8276, B2 => 
                           n10479, ZN => n2299);
   U10415 : OAI22_X1 port map( A1 => n11353, A2 => n11601, B1 => n8275, B2 => 
                           n10479, ZN => n2300);
   U10416 : OAI22_X1 port map( A1 => n11353, A2 => n11609, B1 => n8274, B2 => 
                           n10479, ZN => n2301);
   U10417 : NOR3_X1 port map( A1 => n8273, A2 => Addr_RD2(1), A3 => n8271, ZN 
                           => n10473);
   U10418 : NOR3_X1 port map( A1 => n8269, A2 => Addr_RD1(1), A3 => n8267, ZN 
                           => n9883);
   U10419 : NOR2_X1 port map( A1 => Addr_RD2(4), A2 => Addr_RD2(3), ZN => 
                           n10472);
   U10420 : NOR2_X1 port map( A1 => Addr_RD1(4), A2 => Addr_RD1(3), ZN => n9882
                           );
   U10421 : NOR2_X1 port map( A1 => n8270, A2 => Addr_RD2(4), ZN => n10474);
   U10422 : NOR2_X1 port map( A1 => n8266, A2 => Addr_RD1(4), ZN => n9884);
   U10423 : NOR3_X1 port map( A1 => Addr_RD2(0), A2 => Addr_RD2(2), A3 => n8272
                           , ZN => n10463);
   U10424 : NOR3_X1 port map( A1 => Addr_RD1(0), A2 => Addr_RD1(2), A3 => n8268
                           , ZN => n9873);
   U10425 : NOR3_X1 port map( A1 => Addr_RD2(0), A2 => Addr_RD2(1), A3 => n8271
                           , ZN => n10460);
   U10426 : NOR3_X1 port map( A1 => Addr_RD1(0), A2 => Addr_RD1(1), A3 => n8267
                           , ZN => n9870);
   U10427 : NOR3_X1 port map( A1 => n8273, A2 => Addr_RD2(2), A3 => n8272, ZN 
                           => n10456);
   U10428 : NOR3_X1 port map( A1 => n8269, A2 => Addr_RD1(2), A3 => n8268, ZN 
                           => n9866);
   U10429 : NOR3_X1 port map( A1 => Addr_RD2(1), A2 => Addr_RD2(2), A3 => n8273
                           , ZN => n10454);
   U10430 : NOR3_X1 port map( A1 => Addr_RD1(1), A2 => Addr_RD1(2), A3 => n8269
                           , ZN => n9864);
   U10431 : NOR3_X1 port map( A1 => n8272, A2 => Addr_RD2(0), A3 => n8271, ZN 
                           => n10461);
   U10432 : NOR3_X1 port map( A1 => Addr_RD2(1), A2 => Addr_RD2(2), A3 => 
                           Addr_RD2(0), ZN => n10464);
   U10433 : NOR3_X1 port map( A1 => n8268, A2 => Addr_RD1(0), A3 => n8267, ZN 
                           => n9871);
   U10434 : NOR3_X1 port map( A1 => Addr_RD1(1), A2 => Addr_RD1(2), A3 => 
                           Addr_RD1(0), ZN => n9874);
   U10435 : NAND2_X1 port map( A1 => Addr_WR(1), A2 => Addr_WR(0), ZN => n10518
                           );
   U10436 : NAND2_X1 port map( A1 => Addr_WR(1), A2 => n8265, ZN => n10516);
   U10437 : NAND2_X1 port map( A1 => Addr_WR(0), A2 => n8264, ZN => n10514);
   U10438 : AND2_X1 port map( A1 => Addr_RD2(4), A2 => n8270, ZN => n10457);
   U10439 : AND2_X1 port map( A1 => Addr_RD1(4), A2 => n8266, ZN => n9867);
   U10440 : AND2_X1 port map( A1 => Addr_RD2(4), A2 => Addr_RD2(3), ZN => 
                           n10455);
   U10441 : AND2_X1 port map( A1 => Addr_RD1(4), A2 => Addr_RD1(3), ZN => n9865
                           );
   U10442 : INV_X1 port map( A => Addr_RD2(2), ZN => n8271);
   U10443 : INV_X1 port map( A => Addr_RD1(2), ZN => n8267);
   U10444 : INV_X1 port map( A => Addr_RD2(1), ZN => n8272);
   U10445 : INV_X1 port map( A => Addr_RD1(1), ZN => n8268);
   U10446 : INV_X1 port map( A => Addr_RD2(0), ZN => n8273);
   U10447 : INV_X1 port map( A => Addr_RD1(0), ZN => n8269);
   U10448 : AND3_X1 port map( A1 => WR, A2 => En, A3 => Addr_WR(4), ZN => 
                           n10540);
   U10449 : AND3_X1 port map( A1 => En, A2 => n8261, A3 => WR, ZN => n10519);
   U10450 : INV_X1 port map( A => Addr_WR(4), ZN => n8261);
   U10451 : INV_X1 port map( A => Addr_WR(3), ZN => n8262);
   U10452 : INV_X1 port map( A => Addr_WR(2), ZN => n8263);
   U10453 : INV_X1 port map( A => Addr_WR(0), ZN => n8265);
   U10454 : AOI21_X1 port map( B1 => RD2, B2 => En, A => Rst, ZN => n9909);
   U10455 : AOI21_X1 port map( B1 => RD1, B2 => En, A => Rst, ZN => n9319);
   U10456 : INV_X1 port map( A => Addr_WR(1), ZN => n8264);
   U10457 : NAND2_X1 port map( A1 => DataIN(0), A2 => n11892, ZN => n10510);
   U10458 : NAND2_X1 port map( A1 => DataIN(1), A2 => n11892, ZN => n10509);
   U10459 : NAND2_X1 port map( A1 => DataIN(2), A2 => n11892, ZN => n10508);
   U10460 : NAND2_X1 port map( A1 => DataIN(3), A2 => n11892, ZN => n10507);
   U10461 : NAND2_X1 port map( A1 => DataIN(4), A2 => n11892, ZN => n10506);
   U10462 : NAND2_X1 port map( A1 => DataIN(5), A2 => n11892, ZN => n10505);
   U10463 : NAND2_X1 port map( A1 => DataIN(6), A2 => n11892, ZN => n10504);
   U10464 : NAND2_X1 port map( A1 => DataIN(7), A2 => n11892, ZN => n10503);
   U10465 : NAND2_X1 port map( A1 => DataIN(8), A2 => n11891, ZN => n10502);
   U10466 : NAND2_X1 port map( A1 => DataIN(9), A2 => n11891, ZN => n10501);
   U10467 : NAND2_X1 port map( A1 => DataIN(10), A2 => n11891, ZN => n10500);
   U10468 : NAND2_X1 port map( A1 => DataIN(11), A2 => n11891, ZN => n10499);
   U10469 : NAND2_X1 port map( A1 => DataIN(12), A2 => n11891, ZN => n10498);
   U10470 : NAND2_X1 port map( A1 => DataIN(13), A2 => n11891, ZN => n10497);
   U10471 : NAND2_X1 port map( A1 => DataIN(14), A2 => n11891, ZN => n10496);
   U10472 : NAND2_X1 port map( A1 => DataIN(15), A2 => n11891, ZN => n10495);
   U10473 : NAND2_X1 port map( A1 => DataIN(16), A2 => n11891, ZN => n10494);
   U10474 : NAND2_X1 port map( A1 => DataIN(17), A2 => n11891, ZN => n10493);
   U10475 : NAND2_X1 port map( A1 => DataIN(18), A2 => n11891, ZN => n10492);
   U10476 : NAND2_X1 port map( A1 => DataIN(19), A2 => n11891, ZN => n10491);
   U10477 : NAND2_X1 port map( A1 => DataIN(20), A2 => n11890, ZN => n10490);
   U10478 : NAND2_X1 port map( A1 => DataIN(21), A2 => n11890, ZN => n10489);
   U10479 : NAND2_X1 port map( A1 => DataIN(22), A2 => n11890, ZN => n10488);
   U10480 : NAND2_X1 port map( A1 => DataIN(23), A2 => n11890, ZN => n10487);
   U10481 : NAND2_X1 port map( A1 => DataIN(24), A2 => n11890, ZN => n10486);
   U10482 : NAND2_X1 port map( A1 => DataIN(25), A2 => n11890, ZN => n10485);
   U10483 : NAND2_X1 port map( A1 => DataIN(26), A2 => n11890, ZN => n10484);
   U10484 : NAND2_X1 port map( A1 => DataIN(27), A2 => n11890, ZN => n10483);
   U10485 : NAND2_X1 port map( A1 => DataIN(28), A2 => n11890, ZN => n10482);
   U10486 : NAND2_X1 port map( A1 => DataIN(29), A2 => n11890, ZN => n10481);
   U10487 : NAND2_X1 port map( A1 => DataIN(30), A2 => n11890, ZN => n10480);
   U10488 : NAND2_X1 port map( A1 => DataIN(31), A2 => n11890, ZN => n10478);
   U10489 : BUF_X1 port map( A => n9907, Z => n11702);
   U10490 : NOR2_X1 port map( A1 => Rst, A2 => n11692, ZN => n9907);
   U10491 : BUF_X1 port map( A => n9317, Z => n11841);
   U10492 : NOR2_X1 port map( A1 => Rst, A2 => n11831, ZN => n9317);
   U10493 : INV_X1 port map( A => Addr_RD2(3), ZN => n8270);
   U10494 : INV_X1 port map( A => Addr_RD1(3), ZN => n8266);
   U10495 : INV_X1 port map( A => Rst, ZN => n8260);

end SYN_ARCHBEH;
